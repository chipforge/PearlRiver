magic
tech scmos
timestamp 1540531789
<< polysilicon >>
rect 147 161 152 168
rect 147 130 152 137
<< metal1 >>
rect 90 178 100 200
rect 200 178 210 200
rect 90 168 145 178
rect 155 168 210 178
rect 90 120 145 130
rect 155 120 210 130
rect 90 100 100 120
rect 200 100 210 120
<< rndiffusion >>
rect 147 144 152 148
<< rpdiffusion >>
rect 147 150 152 154
<< rpoly >>
rect 147 148 152 150
<< polycontact >>
rect 145 168 155 178
rect 145 120 155 130
<< polyndiff >>
rect 147 137 152 144
<< polypdiff >>
rect 147 154 152 161
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
