magic
tech scmos
timestamp 1539784506
<< polysilicon >>
rect 140 155 160 159
rect 140 141 160 145
<< metal1 >>
rect 80 179 100 200
rect 200 179 220 200
rect 80 159 140 179
rect 160 159 220 179
rect 80 121 140 141
rect 160 121 220 141
rect 80 100 100 121
rect 200 100 220 121
<< rndiffusion >>
rect 140 151 160 155
<< rpdiffusion >>
rect 140 145 160 149
<< rpoly >>
rect 140 149 160 151
<< polycontact >>
rect 140 159 160 179
rect 140 121 160 141
use L500_TPAD_blank  L500_TPAD_blank_2 ./Library/magic
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
