magic
tech scmos
timestamp 1534326485
<< metal1 >>
rect 0 15 8 18
rect 2 14 8 15
rect 4 4 8 14
rect 0 0 12 4
<< end >>
