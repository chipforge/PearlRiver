magic
tech scmos
timestamp 1540998258
use L500_HVNFET_W108_L22_params  L500_HVNFET_W108_L22_params_0 ../../Library/magic
timestamp 1540991124
transform 1 0 0 0 1 350
box 0 0 300 300
use L500_HVPFET_W108_L22_params  L500_HVPFET_W108_L22_params_0 ../../Library/magic
timestamp 1540993816
transform 1 0 0 0 1 0
box 0 0 300 300
<< end >>
