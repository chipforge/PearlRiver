magic
tech scmos
timestamp 1538589449
<< metal1 >>
rect 154 223 158 227
rect 346 223 350 227
rect 361 223 404 227
rect 100 219 142 223
rect 150 219 354 223
rect 0 100 100 150
rect 154 211 350 219
rect 154 207 166 211
rect 170 207 174 211
rect 330 207 334 211
rect 338 207 350 211
rect 154 203 350 207
rect 154 47 166 203
rect 170 195 334 203
rect 170 55 174 195
rect 178 191 182 195
rect 186 191 190 195
rect 314 191 318 195
rect 322 191 334 195
rect 178 187 334 191
rect 178 63 182 187
rect 186 179 318 187
rect 186 175 198 179
rect 202 175 206 179
rect 298 175 302 179
rect 306 175 318 179
rect 186 171 318 175
rect 186 79 198 171
rect 202 163 302 171
rect 202 159 214 163
rect 218 159 222 163
rect 282 159 286 163
rect 290 159 302 163
rect 202 155 302 159
rect 202 95 214 155
rect 218 147 286 155
rect 218 143 230 147
rect 234 143 238 147
rect 266 143 270 147
rect 274 143 286 147
rect 218 139 286 143
rect 218 111 230 139
rect 234 111 270 139
rect 274 111 286 139
rect 218 107 286 111
rect 218 103 230 107
rect 234 103 238 107
rect 266 103 270 107
rect 274 103 286 107
rect 218 95 286 103
rect 290 95 302 155
rect 202 91 302 95
rect 202 87 214 91
rect 218 87 222 91
rect 282 87 286 91
rect 290 87 302 91
rect 202 79 302 87
rect 306 79 318 171
rect 186 75 318 79
rect 186 71 198 75
rect 202 71 206 75
rect 298 71 302 75
rect 306 71 318 75
rect 186 63 318 71
rect 322 63 334 187
rect 178 59 334 63
rect 178 55 182 59
rect 186 55 190 59
rect 314 55 318 59
rect 322 55 334 59
rect 170 47 334 55
rect 338 47 350 203
rect 154 43 350 47
rect 154 39 166 43
rect 170 39 174 43
rect 330 39 334 43
rect 338 39 350 43
rect 154 31 350 39
rect 404 100 504 150
rect 150 27 354 31
rect 154 23 158 27
rect 346 23 350 27
<< metal2 >>
rect 154 223 158 227
rect 346 223 350 227
rect 150 219 354 223
rect 154 215 158 219
rect 162 215 166 219
rect 338 215 342 219
rect 346 215 350 219
rect 154 211 350 215
rect 154 39 158 211
rect 162 207 166 211
rect 170 207 174 211
rect 330 207 334 211
rect 338 207 342 211
rect 162 203 342 207
rect 162 47 166 203
rect 170 199 174 203
rect 178 199 182 203
rect 322 199 326 203
rect 330 199 334 203
rect 170 195 334 199
rect 170 55 174 195
rect 178 191 182 195
rect 186 191 190 195
rect 314 191 318 195
rect 322 191 326 195
rect 178 187 326 191
rect 178 63 182 187
rect 186 183 190 187
rect 194 183 198 187
rect 306 183 310 187
rect 314 183 318 187
rect 186 179 318 183
rect 186 71 190 179
rect 194 175 198 179
rect 202 175 206 179
rect 298 175 302 179
rect 306 175 310 179
rect 194 171 310 175
rect 194 79 198 171
rect 202 167 206 171
rect 210 167 214 171
rect 290 167 294 171
rect 298 167 302 171
rect 202 163 302 167
rect 202 87 206 163
rect 210 159 214 163
rect 218 159 222 163
rect 282 159 286 163
rect 290 159 294 163
rect 210 155 294 159
rect 210 95 214 155
rect 218 151 222 155
rect 226 151 230 155
rect 274 151 278 155
rect 282 151 286 155
rect 218 147 286 151
rect 218 103 222 147
rect 226 143 230 147
rect 234 143 238 147
rect 266 143 270 147
rect 274 143 278 147
rect 226 139 278 143
rect 226 111 230 139
rect 234 135 238 139
rect 242 135 246 139
rect 258 135 262 139
rect 266 135 270 139
rect 234 131 270 135
rect 234 119 238 131
rect 242 119 262 131
rect 266 119 270 131
rect 234 115 270 119
rect 234 111 238 115
rect 242 111 246 115
rect 258 111 262 115
rect 266 111 270 115
rect 274 111 278 139
rect 226 107 278 111
rect 226 103 230 107
rect 234 103 238 107
rect 266 103 270 107
rect 274 103 278 107
rect 282 103 286 147
rect 218 99 286 103
rect 218 95 222 99
rect 226 95 230 99
rect 274 95 278 99
rect 282 95 286 99
rect 290 95 294 155
rect 210 91 294 95
rect 210 87 214 91
rect 218 87 222 91
rect 282 87 286 91
rect 290 87 294 91
rect 298 87 302 163
rect 202 83 302 87
rect 202 79 206 83
rect 210 79 214 83
rect 290 79 294 83
rect 298 79 302 83
rect 306 79 310 171
rect 194 75 310 79
rect 194 71 198 75
rect 202 71 206 75
rect 298 71 302 75
rect 306 71 310 75
rect 314 71 318 179
rect 186 67 318 71
rect 186 63 190 67
rect 194 63 198 67
rect 306 63 310 67
rect 314 63 318 67
rect 322 63 326 187
rect 178 59 326 63
rect 178 55 182 59
rect 186 55 190 59
rect 314 55 318 59
rect 322 55 326 59
rect 330 55 334 195
rect 170 51 334 55
rect 170 47 174 51
rect 178 47 182 51
rect 322 47 326 51
rect 330 47 334 51
rect 338 47 342 203
rect 162 43 342 47
rect 162 39 166 43
rect 170 39 174 43
rect 330 39 334 43
rect 338 39 342 43
rect 346 39 350 211
rect 154 35 350 39
rect 154 31 158 35
rect 162 31 166 35
rect 338 31 342 35
rect 346 31 350 35
rect 150 27 354 31
rect 154 23 158 27
rect 346 23 350 27
<< metal3 >>
rect 150 219 354 227
rect 150 215 158 219
rect 162 215 166 219
rect 338 215 342 219
rect 346 215 354 219
rect 150 211 354 215
rect 150 39 158 211
rect 162 203 342 211
rect 162 199 174 203
rect 178 199 182 203
rect 322 199 326 203
rect 330 199 342 203
rect 162 195 342 199
rect 162 55 174 195
rect 178 187 326 195
rect 178 183 190 187
rect 194 183 198 187
rect 306 183 310 187
rect 314 183 326 187
rect 178 179 326 183
rect 178 71 190 179
rect 194 171 310 179
rect 194 167 206 171
rect 210 167 214 171
rect 290 167 294 171
rect 298 167 310 171
rect 194 163 310 167
rect 194 87 206 163
rect 210 155 294 163
rect 210 151 222 155
rect 226 151 230 155
rect 274 151 278 155
rect 282 151 294 155
rect 210 147 294 151
rect 210 103 222 147
rect 226 139 278 147
rect 226 135 238 139
rect 242 135 246 139
rect 258 135 262 139
rect 266 135 278 139
rect 226 131 278 135
rect 226 119 238 131
rect 242 119 262 131
rect 266 119 278 131
rect 226 115 278 119
rect 226 111 238 115
rect 242 111 246 115
rect 258 111 262 115
rect 266 111 278 115
rect 226 103 278 111
rect 282 103 294 147
rect 210 99 294 103
rect 210 95 222 99
rect 226 95 230 99
rect 274 95 278 99
rect 282 95 294 99
rect 210 87 294 95
rect 298 87 310 163
rect 194 83 310 87
rect 194 79 206 83
rect 210 79 214 83
rect 290 79 294 83
rect 298 79 310 83
rect 194 71 310 79
rect 314 71 326 179
rect 178 67 326 71
rect 178 63 190 67
rect 194 63 198 67
rect 306 63 310 67
rect 314 63 326 67
rect 178 55 326 63
rect 330 55 342 195
rect 162 51 342 55
rect 162 47 174 51
rect 178 47 182 51
rect 322 47 326 51
rect 330 47 342 51
rect 162 39 342 47
rect 346 39 354 211
rect 150 35 354 39
rect 150 31 158 35
rect 162 31 166 35
rect 338 31 342 35
rect 346 31 354 35
rect 150 23 354 31
<< rpoly >>
rect 167 224 357 226
rect 146 220 157 222
rect 155 210 157 220
rect 167 214 169 224
rect 175 220 193 222
rect 175 214 177 220
rect 191 214 193 220
rect 207 220 225 222
rect 207 214 209 220
rect 223 214 225 220
rect 239 220 257 222
rect 239 214 241 220
rect 255 214 257 220
rect 271 220 289 222
rect 271 214 273 220
rect 287 214 289 220
rect 303 220 321 222
rect 303 214 305 220
rect 319 214 321 220
rect 335 220 349 222
rect 335 214 337 220
rect 167 212 177 214
rect 183 212 193 214
rect 199 212 209 214
rect 215 212 225 214
rect 231 212 241 214
rect 246 212 257 214
rect 263 212 273 214
rect 279 212 289 214
rect 295 212 305 214
rect 311 212 321 214
rect 327 212 337 214
rect 155 208 165 210
rect 163 202 165 208
rect 163 200 173 202
rect 171 194 173 200
rect 183 198 185 212
rect 199 206 201 212
rect 215 206 217 212
rect 231 206 233 212
rect 246 206 248 212
rect 263 206 265 212
rect 279 206 281 212
rect 295 206 297 212
rect 311 206 313 212
rect 327 206 329 212
rect 347 210 349 220
rect 191 204 201 206
rect 207 204 217 206
rect 223 204 233 206
rect 239 204 248 206
rect 255 204 265 206
rect 271 204 281 206
rect 287 204 297 206
rect 303 204 313 206
rect 319 204 329 206
rect 339 208 349 210
rect 191 198 193 204
rect 207 198 209 204
rect 223 198 225 204
rect 239 198 241 204
rect 255 198 257 204
rect 271 198 273 204
rect 287 198 289 204
rect 303 198 305 204
rect 319 198 321 204
rect 339 202 341 208
rect 339 200 349 202
rect 183 196 193 198
rect 199 196 209 198
rect 215 196 225 198
rect 231 196 241 198
rect 246 196 257 198
rect 263 196 273 198
rect 279 196 289 198
rect 295 196 305 198
rect 311 196 321 198
rect 155 192 165 194
rect 171 192 181 194
rect 155 178 157 192
rect 163 186 165 192
rect 179 186 181 192
rect 163 184 173 186
rect 179 184 189 186
rect 171 178 173 184
rect 187 178 189 184
rect 199 182 201 196
rect 215 190 217 196
rect 231 190 233 196
rect 246 190 248 196
rect 263 190 265 196
rect 279 190 281 196
rect 295 190 297 196
rect 311 190 313 196
rect 207 188 217 190
rect 223 188 233 190
rect 239 188 248 190
rect 255 188 265 190
rect 271 188 281 190
rect 287 188 297 190
rect 303 188 313 190
rect 323 192 341 194
rect 207 182 209 188
rect 223 182 225 188
rect 239 182 241 188
rect 255 182 257 188
rect 271 182 273 188
rect 287 182 289 188
rect 303 182 305 188
rect 323 186 325 192
rect 339 186 341 192
rect 347 186 349 200
rect 323 184 333 186
rect 339 184 349 186
rect 199 180 209 182
rect 215 180 225 182
rect 231 180 241 182
rect 246 180 257 182
rect 263 180 273 182
rect 279 180 289 182
rect 295 180 305 182
rect 155 176 165 178
rect 171 176 181 178
rect 187 176 197 178
rect 163 170 165 176
rect 179 170 181 176
rect 195 170 197 176
rect 163 168 173 170
rect 179 168 189 170
rect 195 168 205 170
rect 171 162 173 168
rect 187 162 189 168
rect 203 162 205 168
rect 215 166 217 180
rect 231 174 233 180
rect 246 174 248 180
rect 263 174 265 180
rect 279 174 281 180
rect 295 174 297 180
rect 331 178 333 184
rect 223 172 233 174
rect 239 172 248 174
rect 255 172 265 174
rect 271 172 281 174
rect 287 172 297 174
rect 307 176 325 178
rect 331 176 341 178
rect 223 166 225 172
rect 239 166 241 172
rect 255 166 257 172
rect 271 166 273 172
rect 287 166 289 172
rect 307 170 309 176
rect 323 170 325 176
rect 339 170 341 176
rect 307 168 317 170
rect 323 168 333 170
rect 339 168 349 170
rect 215 164 225 166
rect 231 164 241 166
rect 246 164 257 166
rect 263 164 273 166
rect 279 164 289 166
rect 155 160 165 162
rect 171 160 181 162
rect 187 160 197 162
rect 203 160 213 162
rect 155 146 157 160
rect 163 154 165 160
rect 179 154 181 160
rect 195 154 197 160
rect 211 154 213 160
rect 163 152 173 154
rect 179 152 189 154
rect 195 152 205 154
rect 211 152 221 154
rect 171 146 173 152
rect 187 146 189 152
rect 203 146 205 152
rect 219 146 221 152
rect 231 150 233 164
rect 246 158 248 164
rect 263 158 265 164
rect 279 158 281 164
rect 315 162 317 168
rect 331 162 333 168
rect 239 156 248 158
rect 255 156 265 158
rect 271 156 281 158
rect 291 160 309 162
rect 315 160 325 162
rect 331 160 341 162
rect 239 150 241 156
rect 255 150 257 156
rect 271 150 273 156
rect 291 154 293 160
rect 307 154 309 160
rect 323 154 325 160
rect 339 154 341 160
rect 347 154 349 168
rect 291 152 301 154
rect 307 152 317 154
rect 323 152 333 154
rect 339 152 349 154
rect 231 148 241 150
rect 247 148 257 150
rect 263 148 273 150
rect 155 144 165 146
rect 171 144 181 146
rect 187 144 197 146
rect 203 144 213 146
rect 219 144 229 146
rect 163 138 165 144
rect 179 138 181 144
rect 195 138 197 144
rect 211 138 213 144
rect 227 138 229 144
rect 163 136 173 138
rect 179 136 189 138
rect 195 136 205 138
rect 211 136 221 138
rect 227 136 237 138
rect 171 130 173 136
rect 187 130 189 136
rect 203 130 205 136
rect 219 130 221 136
rect 235 130 237 136
rect 247 134 249 148
rect 263 142 265 148
rect 299 146 301 152
rect 315 146 317 152
rect 331 146 333 152
rect 255 140 265 142
rect 275 144 293 146
rect 299 144 309 146
rect 315 144 325 146
rect 331 144 341 146
rect 255 134 257 140
rect 275 138 277 144
rect 291 138 293 144
rect 307 138 309 144
rect 323 138 325 144
rect 339 138 341 144
rect 275 136 285 138
rect 291 136 301 138
rect 307 136 317 138
rect 323 136 333 138
rect 339 136 349 138
rect 247 132 257 134
rect 283 130 285 136
rect 299 130 301 136
rect 315 130 317 136
rect 331 130 333 136
rect 155 128 165 130
rect 171 128 181 130
rect 187 128 197 130
rect 203 128 213 130
rect 219 128 229 130
rect 235 128 245 130
rect 155 114 157 128
rect 163 122 165 128
rect 179 122 181 128
rect 195 122 197 128
rect 211 122 213 128
rect 227 122 229 128
rect 243 122 245 128
rect 163 120 173 122
rect 179 120 189 122
rect 195 120 205 122
rect 211 120 221 122
rect 227 120 245 122
rect 259 128 277 130
rect 283 128 293 130
rect 299 128 309 130
rect 315 128 325 130
rect 331 128 341 130
rect 259 122 261 128
rect 275 122 277 128
rect 291 122 293 128
rect 307 122 309 128
rect 323 122 325 128
rect 339 122 341 128
rect 347 122 349 136
rect 259 120 269 122
rect 275 120 285 122
rect 291 120 301 122
rect 307 120 317 122
rect 323 120 333 122
rect 339 120 349 122
rect 171 114 173 120
rect 187 114 189 120
rect 203 114 205 120
rect 219 114 221 120
rect 247 116 257 118
rect 155 112 165 114
rect 171 112 181 114
rect 187 112 197 114
rect 203 112 213 114
rect 219 112 229 114
rect 163 106 165 112
rect 179 106 181 112
rect 195 106 197 112
rect 211 106 213 112
rect 227 106 229 112
rect 247 110 249 116
rect 163 104 173 106
rect 179 104 189 106
rect 195 104 205 106
rect 211 104 229 106
rect 239 108 249 110
rect 171 98 173 104
rect 187 98 189 104
rect 203 98 205 104
rect 239 102 241 108
rect 255 102 257 116
rect 267 114 269 120
rect 283 114 285 120
rect 299 114 301 120
rect 315 114 317 120
rect 331 114 333 120
rect 267 112 277 114
rect 283 112 293 114
rect 299 112 309 114
rect 315 112 325 114
rect 331 112 341 114
rect 275 106 277 112
rect 291 106 293 112
rect 307 106 309 112
rect 323 106 325 112
rect 339 106 341 112
rect 275 104 285 106
rect 291 104 301 106
rect 307 104 317 106
rect 323 104 333 106
rect 339 104 349 106
rect 231 100 241 102
rect 247 100 257 102
rect 263 100 273 102
rect 155 96 165 98
rect 171 96 181 98
rect 187 96 197 98
rect 203 96 213 98
rect 155 82 157 96
rect 163 90 165 96
rect 179 90 181 96
rect 195 90 197 96
rect 211 90 213 96
rect 231 94 233 100
rect 247 94 249 100
rect 263 94 265 100
rect 163 88 173 90
rect 179 88 189 90
rect 195 88 213 90
rect 223 92 233 94
rect 239 92 249 94
rect 255 92 265 94
rect 171 82 173 88
rect 187 82 189 88
rect 223 86 225 92
rect 239 86 241 92
rect 255 86 257 92
rect 271 86 273 100
rect 283 98 285 104
rect 299 98 301 104
rect 315 98 317 104
rect 331 98 333 104
rect 283 96 293 98
rect 299 96 309 98
rect 315 96 325 98
rect 331 96 341 98
rect 291 90 293 96
rect 307 90 309 96
rect 323 90 325 96
rect 339 90 341 96
rect 347 90 349 104
rect 291 88 301 90
rect 307 88 317 90
rect 323 88 333 90
rect 339 88 349 90
rect 215 84 225 86
rect 231 84 241 86
rect 247 84 257 86
rect 263 84 273 86
rect 279 84 289 86
rect 155 80 165 82
rect 171 80 181 82
rect 187 80 197 82
rect 163 74 165 80
rect 179 74 181 80
rect 195 74 197 80
rect 215 78 217 84
rect 231 78 233 84
rect 247 78 249 84
rect 263 78 265 84
rect 279 78 281 84
rect 163 72 173 74
rect 179 72 197 74
rect 207 76 217 78
rect 223 76 233 78
rect 239 76 249 78
rect 255 76 265 78
rect 271 76 281 78
rect 171 66 173 72
rect 207 70 209 76
rect 223 70 225 76
rect 239 70 241 76
rect 255 70 257 76
rect 271 70 273 76
rect 287 70 289 84
rect 299 82 301 88
rect 315 82 317 88
rect 331 82 333 88
rect 299 80 309 82
rect 315 80 325 82
rect 331 80 341 82
rect 307 74 309 80
rect 323 74 325 80
rect 339 74 341 80
rect 307 72 317 74
rect 323 72 333 74
rect 339 72 349 74
rect 199 68 209 70
rect 215 68 225 70
rect 231 68 241 70
rect 247 68 257 70
rect 263 68 273 70
rect 279 68 289 70
rect 295 68 305 70
rect 155 64 165 66
rect 171 64 181 66
rect 155 50 157 64
rect 163 58 165 64
rect 179 58 181 64
rect 199 62 201 68
rect 215 62 217 68
rect 231 62 233 68
rect 247 62 249 68
rect 263 62 265 68
rect 279 62 281 68
rect 295 62 297 68
rect 163 56 181 58
rect 191 60 201 62
rect 207 60 217 62
rect 223 60 233 62
rect 239 60 249 62
rect 255 60 265 62
rect 271 60 281 62
rect 287 60 297 62
rect 191 54 193 60
rect 207 54 209 60
rect 223 54 225 60
rect 239 54 241 60
rect 255 54 257 60
rect 271 54 273 60
rect 287 54 289 60
rect 303 54 305 68
rect 315 66 317 72
rect 331 66 333 72
rect 315 64 325 66
rect 331 64 341 66
rect 323 58 325 64
rect 339 58 341 64
rect 347 58 349 72
rect 323 56 333 58
rect 339 56 349 58
rect 183 52 193 54
rect 199 52 209 54
rect 215 52 225 54
rect 231 52 241 54
rect 247 52 257 54
rect 263 52 273 54
rect 279 52 289 54
rect 295 52 305 54
rect 311 52 321 54
rect 155 48 165 50
rect 163 42 165 48
rect 183 46 185 52
rect 199 46 201 52
rect 215 46 217 52
rect 231 46 233 52
rect 247 46 249 52
rect 263 46 265 52
rect 279 46 281 52
rect 295 46 297 52
rect 311 46 313 52
rect 155 40 165 42
rect 175 44 185 46
rect 191 44 201 46
rect 207 44 217 46
rect 223 44 233 46
rect 239 44 249 46
rect 255 44 265 46
rect 271 44 281 46
rect 287 44 297 46
rect 303 44 313 46
rect 155 30 157 40
rect 175 38 177 44
rect 191 38 193 44
rect 207 38 209 44
rect 223 38 225 44
rect 239 38 241 44
rect 255 38 257 44
rect 271 38 273 44
rect 287 38 289 44
rect 303 38 305 44
rect 319 38 321 52
rect 331 50 333 56
rect 331 48 341 50
rect 339 42 341 48
rect 339 40 349 42
rect 167 36 177 38
rect 183 36 193 38
rect 199 36 209 38
rect 215 36 225 38
rect 232 36 241 38
rect 247 36 257 38
rect 263 36 273 38
rect 279 36 289 38
rect 296 36 305 38
rect 311 36 321 38
rect 327 36 337 38
rect 167 30 169 36
rect 155 28 169 30
rect 183 30 185 36
rect 199 30 201 36
rect 183 28 201 30
rect 215 30 217 36
rect 232 30 234 36
rect 215 28 234 30
rect 247 30 249 36
rect 263 30 265 36
rect 247 28 265 30
rect 279 30 281 36
rect 296 30 298 36
rect 279 28 298 30
rect 311 30 313 36
rect 327 30 329 36
rect 311 28 329 30
rect 335 30 337 36
rect 347 30 349 40
rect 335 28 349 30
<< polycontact >>
rect 142 219 146 223
rect 357 223 361 227
<< m2contact >>
rect 150 223 154 227
rect 158 223 346 227
rect 350 223 354 227
rect 150 31 154 219
rect 166 207 170 211
rect 174 207 330 211
rect 334 207 338 211
rect 166 47 170 203
rect 182 191 186 195
rect 190 191 314 195
rect 318 191 322 195
rect 182 63 186 187
rect 198 175 202 179
rect 206 175 298 179
rect 302 175 306 179
rect 198 79 202 171
rect 214 159 218 163
rect 222 159 282 163
rect 286 159 290 163
rect 214 95 218 155
rect 230 143 234 147
rect 238 143 266 147
rect 270 143 274 147
rect 230 111 234 139
rect 270 111 274 139
rect 230 103 234 107
rect 238 103 266 107
rect 270 103 274 107
rect 286 95 290 155
rect 214 87 218 91
rect 222 87 282 91
rect 286 87 290 91
rect 302 79 306 171
rect 198 71 202 75
rect 206 71 298 75
rect 302 71 306 75
rect 318 63 322 187
rect 182 55 186 59
rect 190 55 314 59
rect 318 55 322 59
rect 334 47 338 203
rect 166 39 170 43
rect 174 39 330 43
rect 334 39 338 43
rect 350 31 354 219
rect 150 23 154 27
rect 158 23 346 27
rect 350 23 354 27
<< m3contact >>
rect 158 215 162 219
rect 166 215 338 219
rect 342 215 346 219
rect 158 39 162 211
rect 174 199 178 203
rect 182 199 322 203
rect 326 199 330 203
rect 174 55 178 195
rect 190 183 194 187
rect 198 183 306 187
rect 310 183 314 187
rect 190 71 194 179
rect 206 167 210 171
rect 214 167 290 171
rect 294 167 298 171
rect 206 87 210 163
rect 222 151 226 155
rect 230 151 274 155
rect 278 151 282 155
rect 222 103 226 147
rect 238 135 242 139
rect 246 135 258 139
rect 262 135 266 139
rect 238 119 242 131
rect 262 119 266 131
rect 238 111 242 115
rect 246 111 258 115
rect 262 111 266 115
rect 278 103 282 147
rect 222 95 226 99
rect 230 95 274 99
rect 278 95 282 99
rect 294 87 298 163
rect 206 79 210 83
rect 214 79 290 83
rect 294 79 298 83
rect 310 71 314 179
rect 190 63 194 67
rect 198 63 306 67
rect 310 63 314 67
rect 326 55 330 195
rect 174 47 178 51
rect 182 47 322 51
rect 326 47 330 51
rect 342 39 346 211
rect 158 31 162 35
rect 166 31 338 35
rect 342 31 346 35
<< glass >>
rect 162 35 342 215
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 0 0 1 150
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 404 0 1 150
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 404 0 1 0
box 0 0 100 100
<< end >>
