magic
tech scmos
timestamp 1533657739
<< metal3 >>
rect 90 117 91 118
rect 91 117 92 118
rect 92 117 93 118
rect 89 116 90 117
rect 90 116 91 117
rect 91 116 92 117
rect 92 116 93 117
rect 88 115 89 116
rect 89 115 90 116
rect 90 115 91 116
rect 91 115 92 116
rect 92 115 93 116
rect 93 115 94 116
rect 88 114 89 115
rect 89 114 90 115
rect 90 114 91 115
rect 91 114 92 115
rect 92 114 93 115
rect 93 114 94 115
rect 87 113 88 114
rect 88 113 89 114
rect 89 113 90 114
rect 90 113 91 114
rect 91 113 92 114
rect 92 113 93 114
rect 93 113 94 114
rect 94 113 95 114
rect 86 112 87 113
rect 87 112 88 113
rect 88 112 89 113
rect 89 112 90 113
rect 90 112 91 113
rect 91 112 92 113
rect 92 112 93 113
rect 93 112 94 113
rect 94 112 95 113
rect 86 111 87 112
rect 87 111 88 112
rect 88 111 89 112
rect 89 111 90 112
rect 90 111 91 112
rect 91 111 92 112
rect 92 111 93 112
rect 93 111 94 112
rect 94 111 95 112
rect 84 110 85 111
rect 85 110 86 111
rect 86 110 87 111
rect 87 110 88 111
rect 88 110 89 111
rect 89 110 90 111
rect 90 110 91 111
rect 91 110 92 111
rect 92 110 93 111
rect 93 110 94 111
rect 94 110 95 111
rect 54 109 55 110
rect 55 109 56 110
rect 56 109 57 110
rect 57 109 58 110
rect 58 109 59 110
rect 59 109 60 110
rect 60 109 61 110
rect 61 109 62 110
rect 62 109 63 110
rect 63 109 64 110
rect 64 109 65 110
rect 84 109 85 110
rect 85 109 86 110
rect 86 109 87 110
rect 87 109 88 110
rect 88 109 89 110
rect 89 109 90 110
rect 90 109 91 110
rect 91 109 92 110
rect 92 109 93 110
rect 93 109 94 110
rect 94 109 95 110
rect 52 108 53 109
rect 53 108 54 109
rect 54 108 55 109
rect 55 108 56 109
rect 56 108 57 109
rect 57 108 58 109
rect 58 108 59 109
rect 59 108 60 109
rect 60 108 61 109
rect 61 108 62 109
rect 62 108 63 109
rect 63 108 64 109
rect 64 108 65 109
rect 65 108 66 109
rect 66 108 67 109
rect 67 108 68 109
rect 68 108 69 109
rect 83 108 84 109
rect 84 108 85 109
rect 85 108 86 109
rect 86 108 87 109
rect 87 108 88 109
rect 88 108 89 109
rect 89 108 90 109
rect 90 108 91 109
rect 91 108 92 109
rect 92 108 93 109
rect 93 108 94 109
rect 94 108 95 109
rect 50 107 51 108
rect 51 107 52 108
rect 52 107 53 108
rect 53 107 54 108
rect 54 107 55 108
rect 55 107 56 108
rect 56 107 57 108
rect 57 107 58 108
rect 58 107 59 108
rect 59 107 60 108
rect 60 107 61 108
rect 62 107 63 108
rect 63 107 64 108
rect 64 107 65 108
rect 65 107 66 108
rect 66 107 67 108
rect 67 107 68 108
rect 68 107 69 108
rect 69 107 70 108
rect 70 107 71 108
rect 82 107 83 108
rect 83 107 84 108
rect 84 107 85 108
rect 85 107 86 108
rect 86 107 87 108
rect 87 107 88 108
rect 88 107 89 108
rect 89 107 90 108
rect 90 107 91 108
rect 91 107 92 108
rect 92 107 93 108
rect 93 107 94 108
rect 94 107 95 108
rect 49 106 50 107
rect 50 106 51 107
rect 51 106 52 107
rect 68 106 69 107
rect 69 106 70 107
rect 70 106 71 107
rect 71 106 72 107
rect 72 106 73 107
rect 81 106 82 107
rect 82 106 83 107
rect 83 106 84 107
rect 84 106 85 107
rect 85 106 86 107
rect 88 106 89 107
rect 89 106 90 107
rect 90 106 91 107
rect 91 106 92 107
rect 92 106 93 107
rect 93 106 94 107
rect 94 106 95 107
rect 49 105 50 106
rect 69 105 70 106
rect 70 105 71 106
rect 71 105 72 106
rect 72 105 73 106
rect 73 105 74 106
rect 80 105 81 106
rect 81 105 82 106
rect 82 105 83 106
rect 83 105 84 106
rect 84 105 85 106
rect 88 105 89 106
rect 89 105 90 106
rect 90 105 91 106
rect 91 105 92 106
rect 92 105 93 106
rect 93 105 94 106
rect 94 105 95 106
rect 47 104 48 105
rect 70 104 71 105
rect 71 104 72 105
rect 72 104 73 105
rect 73 104 74 105
rect 74 104 75 105
rect 80 104 81 105
rect 81 104 82 105
rect 82 104 83 105
rect 83 104 84 105
rect 88 104 89 105
rect 89 104 90 105
rect 90 104 91 105
rect 91 104 92 105
rect 92 104 93 105
rect 93 104 94 105
rect 94 104 95 105
rect 45 103 46 104
rect 46 103 47 104
rect 47 103 48 104
rect 72 103 73 104
rect 73 103 74 104
rect 74 103 75 104
rect 75 103 76 104
rect 78 103 79 104
rect 79 103 80 104
rect 80 103 81 104
rect 81 103 82 104
rect 82 103 83 104
rect 88 103 89 104
rect 89 103 90 104
rect 90 103 91 104
rect 91 103 92 104
rect 92 103 93 104
rect 93 103 94 104
rect 94 103 95 104
rect 45 102 46 103
rect 46 102 47 103
rect 73 102 74 103
rect 74 102 75 103
rect 75 102 76 103
rect 76 102 77 103
rect 77 102 78 103
rect 78 102 79 103
rect 79 102 80 103
rect 80 102 81 103
rect 81 102 82 103
rect 88 102 89 103
rect 89 102 90 103
rect 90 102 91 103
rect 91 102 92 103
rect 92 102 93 103
rect 93 102 94 103
rect 94 102 95 103
rect 44 101 45 102
rect 45 101 46 102
rect 74 101 75 102
rect 75 101 76 102
rect 76 101 77 102
rect 77 101 78 102
rect 78 101 79 102
rect 79 101 80 102
rect 80 101 81 102
rect 81 101 82 102
rect 87 101 88 102
rect 88 101 89 102
rect 89 101 90 102
rect 90 101 91 102
rect 91 101 92 102
rect 92 101 93 102
rect 42 100 43 101
rect 43 100 44 101
rect 44 100 45 101
rect 74 100 75 101
rect 75 100 76 101
rect 76 100 77 101
rect 77 100 78 101
rect 78 100 79 101
rect 79 100 80 101
rect 80 100 81 101
rect 87 100 88 101
rect 88 100 89 101
rect 89 100 90 101
rect 90 100 91 101
rect 41 99 42 100
rect 42 99 43 100
rect 43 99 44 100
rect 74 99 75 100
rect 75 99 76 100
rect 76 99 77 100
rect 77 99 78 100
rect 78 99 79 100
rect 79 99 80 100
rect 86 99 87 100
rect 87 99 88 100
rect 88 99 89 100
rect 41 98 42 99
rect 42 98 43 99
rect 43 98 44 99
rect 73 98 74 99
rect 74 98 75 99
rect 75 98 76 99
rect 76 98 77 99
rect 77 98 78 99
rect 78 98 79 99
rect 79 98 80 99
rect 85 98 86 99
rect 86 98 87 99
rect 87 98 88 99
rect 39 97 40 98
rect 40 97 41 98
rect 41 97 42 98
rect 73 97 74 98
rect 74 97 75 98
rect 75 97 76 98
rect 76 97 77 98
rect 77 97 78 98
rect 78 97 79 98
rect 83 97 84 98
rect 84 97 85 98
rect 85 97 86 98
rect 86 97 87 98
rect 39 96 40 97
rect 40 96 41 97
rect 73 96 74 97
rect 74 96 75 97
rect 75 96 76 97
rect 76 96 77 97
rect 77 96 78 97
rect 82 96 83 97
rect 83 96 84 97
rect 84 96 85 97
rect 85 96 86 97
rect 38 95 39 96
rect 39 95 40 96
rect 73 95 74 96
rect 74 95 75 96
rect 75 95 76 96
rect 76 95 77 96
rect 77 95 78 96
rect 81 95 82 96
rect 82 95 83 96
rect 83 95 84 96
rect 84 95 85 96
rect 36 94 37 95
rect 37 94 38 95
rect 38 94 39 95
rect 39 94 40 95
rect 72 94 73 95
rect 73 94 74 95
rect 74 94 75 95
rect 75 94 76 95
rect 76 94 77 95
rect 79 94 80 95
rect 80 94 81 95
rect 81 94 82 95
rect 82 94 83 95
rect 83 94 84 95
rect 35 93 36 94
rect 36 93 37 94
rect 37 93 38 94
rect 73 93 74 94
rect 74 93 75 94
rect 75 93 76 94
rect 76 93 77 94
rect 78 93 79 94
rect 79 93 80 94
rect 80 93 81 94
rect 81 93 82 94
rect 82 93 83 94
rect 34 92 35 93
rect 35 92 36 93
rect 36 92 37 93
rect 72 92 73 93
rect 73 92 74 93
rect 74 92 75 93
rect 75 92 76 93
rect 76 92 77 93
rect 78 92 79 93
rect 79 92 80 93
rect 80 92 81 93
rect 81 92 82 93
rect 33 91 34 92
rect 34 91 35 92
rect 35 91 36 92
rect 47 91 48 92
rect 48 91 49 92
rect 49 91 50 92
rect 50 91 51 92
rect 51 91 52 92
rect 52 91 53 92
rect 53 91 54 92
rect 54 91 55 92
rect 55 91 56 92
rect 72 91 73 92
rect 73 91 74 92
rect 74 91 75 92
rect 75 91 76 92
rect 76 91 77 92
rect 77 91 78 92
rect 78 91 79 92
rect 79 91 80 92
rect 80 91 81 92
rect 32 90 33 91
rect 33 90 34 91
rect 34 90 35 91
rect 45 90 46 91
rect 46 90 47 91
rect 47 90 48 91
rect 48 90 49 91
rect 49 90 50 91
rect 50 90 51 91
rect 51 90 52 91
rect 52 90 53 91
rect 53 90 54 91
rect 54 90 55 91
rect 55 90 56 91
rect 56 90 57 91
rect 57 90 58 91
rect 58 90 59 91
rect 59 90 60 91
rect 60 90 61 91
rect 72 90 73 91
rect 73 90 74 91
rect 74 90 75 91
rect 75 90 76 91
rect 76 90 77 91
rect 77 90 78 91
rect 78 90 79 91
rect 79 90 80 91
rect 80 90 81 91
rect 30 89 31 90
rect 31 89 32 90
rect 32 89 33 90
rect 42 89 43 90
rect 43 89 44 90
rect 55 89 56 90
rect 56 89 57 90
rect 57 89 58 90
rect 58 89 59 90
rect 59 89 60 90
rect 60 89 61 90
rect 61 89 62 90
rect 62 89 63 90
rect 72 89 73 90
rect 73 89 74 90
rect 74 89 75 90
rect 75 89 76 90
rect 76 89 77 90
rect 77 89 78 90
rect 78 89 79 90
rect 79 89 80 90
rect 29 88 30 89
rect 30 88 31 89
rect 31 88 32 89
rect 41 88 42 89
rect 42 88 43 89
rect 43 88 44 89
rect 58 88 59 89
rect 59 88 60 89
rect 60 88 61 89
rect 61 88 62 89
rect 62 88 63 89
rect 63 88 64 89
rect 64 88 65 89
rect 72 88 73 89
rect 73 88 74 89
rect 74 88 75 89
rect 75 88 76 89
rect 76 88 77 89
rect 77 88 78 89
rect 78 88 79 89
rect 79 88 80 89
rect 27 87 28 88
rect 28 87 29 88
rect 29 87 30 88
rect 30 87 31 88
rect 39 87 40 88
rect 40 87 41 88
rect 41 87 42 88
rect 42 87 43 88
rect 62 87 63 88
rect 63 87 64 88
rect 64 87 65 88
rect 65 87 66 88
rect 66 87 67 88
rect 67 87 68 88
rect 68 87 69 88
rect 72 87 73 88
rect 73 87 74 88
rect 74 87 75 88
rect 75 87 76 88
rect 76 87 77 88
rect 77 87 78 88
rect 78 87 79 88
rect 26 86 27 87
rect 27 86 28 87
rect 28 86 29 87
rect 29 86 30 87
rect 37 86 38 87
rect 38 86 39 87
rect 39 86 40 87
rect 40 86 41 87
rect 41 86 42 87
rect 66 86 67 87
rect 67 86 68 87
rect 68 86 69 87
rect 69 86 70 87
rect 72 86 73 87
rect 73 86 74 87
rect 74 86 75 87
rect 75 86 76 87
rect 76 86 77 87
rect 77 86 78 87
rect 78 86 79 87
rect 84 86 85 87
rect 95 86 96 87
rect 96 86 97 87
rect 97 86 98 87
rect 98 86 99 87
rect 24 85 25 86
rect 25 85 26 86
rect 26 85 27 86
rect 27 85 28 86
rect 37 85 38 86
rect 38 85 39 86
rect 39 85 40 86
rect 40 85 41 86
rect 69 85 70 86
rect 72 85 73 86
rect 73 85 74 86
rect 74 85 75 86
rect 75 85 76 86
rect 76 85 77 86
rect 77 85 78 86
rect 78 85 79 86
rect 82 85 83 86
rect 83 85 84 86
rect 84 85 85 86
rect 85 85 86 86
rect 86 85 87 86
rect 87 85 88 86
rect 88 85 89 86
rect 89 85 90 86
rect 90 85 91 86
rect 91 85 92 86
rect 92 85 93 86
rect 93 85 94 86
rect 94 85 95 86
rect 95 85 96 86
rect 96 85 97 86
rect 97 85 98 86
rect 98 85 99 86
rect 99 85 100 86
rect 100 85 101 86
rect 101 85 102 86
rect 102 85 103 86
rect 103 85 104 86
rect 104 85 105 86
rect 22 84 23 85
rect 23 84 24 85
rect 24 84 25 85
rect 25 84 26 85
rect 26 84 27 85
rect 35 84 36 85
rect 36 84 37 85
rect 37 84 38 85
rect 38 84 39 85
rect 39 84 40 85
rect 72 84 73 85
rect 73 84 74 85
rect 74 84 75 85
rect 75 84 76 85
rect 76 84 77 85
rect 77 84 78 85
rect 78 84 79 85
rect 80 84 81 85
rect 81 84 82 85
rect 82 84 83 85
rect 83 84 84 85
rect 84 84 85 85
rect 85 84 86 85
rect 86 84 87 85
rect 87 84 88 85
rect 88 84 89 85
rect 89 84 90 85
rect 90 84 91 85
rect 91 84 92 85
rect 92 84 93 85
rect 93 84 94 85
rect 94 84 95 85
rect 95 84 96 85
rect 96 84 97 85
rect 97 84 98 85
rect 98 84 99 85
rect 99 84 100 85
rect 100 84 101 85
rect 101 84 102 85
rect 102 84 103 85
rect 103 84 104 85
rect 104 84 105 85
rect 105 84 106 85
rect 106 84 107 85
rect 107 84 108 85
rect 21 83 22 84
rect 22 83 23 84
rect 23 83 24 84
rect 24 83 25 84
rect 25 83 26 84
rect 34 83 35 84
rect 35 83 36 84
rect 36 83 37 84
rect 37 83 38 84
rect 38 83 39 84
rect 72 83 73 84
rect 73 83 74 84
rect 74 83 75 84
rect 75 83 76 84
rect 76 83 77 84
rect 77 83 78 84
rect 78 83 79 84
rect 79 83 80 84
rect 80 83 81 84
rect 81 83 82 84
rect 82 83 83 84
rect 83 83 84 84
rect 84 83 85 84
rect 85 83 86 84
rect 86 83 87 84
rect 87 83 88 84
rect 88 83 89 84
rect 89 83 90 84
rect 100 83 101 84
rect 101 83 102 84
rect 102 83 103 84
rect 103 83 104 84
rect 104 83 105 84
rect 105 83 106 84
rect 106 83 107 84
rect 107 83 108 84
rect 108 83 109 84
rect 19 82 20 83
rect 20 82 21 83
rect 21 82 22 83
rect 22 82 23 83
rect 23 82 24 83
rect 33 82 34 83
rect 34 82 35 83
rect 35 82 36 83
rect 36 82 37 83
rect 37 82 38 83
rect 72 82 73 83
rect 73 82 74 83
rect 74 82 75 83
rect 75 82 76 83
rect 76 82 77 83
rect 77 82 78 83
rect 78 82 79 83
rect 79 82 80 83
rect 80 82 81 83
rect 81 82 82 83
rect 82 82 83 83
rect 83 82 84 83
rect 84 82 85 83
rect 85 82 86 83
rect 86 82 87 83
rect 102 82 103 83
rect 103 82 104 83
rect 104 82 105 83
rect 105 82 106 83
rect 106 82 107 83
rect 107 82 108 83
rect 108 82 109 83
rect 109 82 110 83
rect 110 82 111 83
rect 17 81 18 82
rect 18 81 19 82
rect 19 81 20 82
rect 20 81 21 82
rect 21 81 22 82
rect 22 81 23 82
rect 32 81 33 82
rect 33 81 34 82
rect 34 81 35 82
rect 35 81 36 82
rect 36 81 37 82
rect 37 81 38 82
rect 72 81 73 82
rect 73 81 74 82
rect 74 81 75 82
rect 75 81 76 82
rect 76 81 77 82
rect 77 81 78 82
rect 78 81 79 82
rect 79 81 80 82
rect 80 81 81 82
rect 81 81 82 82
rect 82 81 83 82
rect 83 81 84 82
rect 84 81 85 82
rect 103 81 104 82
rect 104 81 105 82
rect 105 81 106 82
rect 106 81 107 82
rect 107 81 108 82
rect 108 81 109 82
rect 109 81 110 82
rect 110 81 111 82
rect 14 80 15 81
rect 15 80 16 81
rect 16 80 17 81
rect 17 80 18 81
rect 18 80 19 81
rect 19 80 20 81
rect 20 80 21 81
rect 21 80 22 81
rect 31 80 32 81
rect 32 80 33 81
rect 33 80 34 81
rect 34 80 35 81
rect 35 80 36 81
rect 36 80 37 81
rect 71 80 72 81
rect 72 80 73 81
rect 73 80 74 81
rect 74 80 75 81
rect 75 80 76 81
rect 76 80 77 81
rect 77 80 78 81
rect 78 80 79 81
rect 79 80 80 81
rect 80 80 81 81
rect 81 80 82 81
rect 104 80 105 81
rect 105 80 106 81
rect 106 80 107 81
rect 107 80 108 81
rect 108 80 109 81
rect 109 80 110 81
rect 110 80 111 81
rect 111 80 112 81
rect 13 79 14 80
rect 14 79 15 80
rect 15 79 16 80
rect 16 79 17 80
rect 17 79 18 80
rect 18 79 19 80
rect 30 79 31 80
rect 31 79 32 80
rect 32 79 33 80
rect 33 79 34 80
rect 34 79 35 80
rect 35 79 36 80
rect 70 79 71 80
rect 71 79 72 80
rect 72 79 73 80
rect 73 79 74 80
rect 74 79 75 80
rect 75 79 76 80
rect 76 79 77 80
rect 105 79 106 80
rect 106 79 107 80
rect 107 79 108 80
rect 108 79 109 80
rect 109 79 110 80
rect 110 79 111 80
rect 111 79 112 80
rect 112 79 113 80
rect 11 78 12 79
rect 12 78 13 79
rect 13 78 14 79
rect 14 78 15 79
rect 15 78 16 79
rect 16 78 17 79
rect 17 78 18 79
rect 29 78 30 79
rect 30 78 31 79
rect 31 78 32 79
rect 32 78 33 79
rect 33 78 34 79
rect 34 78 35 79
rect 70 78 71 79
rect 71 78 72 79
rect 72 78 73 79
rect 106 78 107 79
rect 107 78 108 79
rect 108 78 109 79
rect 109 78 110 79
rect 110 78 111 79
rect 111 78 112 79
rect 112 78 113 79
rect 8 77 9 78
rect 9 77 10 78
rect 10 77 11 78
rect 11 77 12 78
rect 12 77 13 78
rect 13 77 14 78
rect 14 77 15 78
rect 15 77 16 78
rect 28 77 29 78
rect 29 77 30 78
rect 30 77 31 78
rect 31 77 32 78
rect 32 77 33 78
rect 33 77 34 78
rect 106 77 107 78
rect 107 77 108 78
rect 108 77 109 78
rect 109 77 110 78
rect 110 77 111 78
rect 111 77 112 78
rect 112 77 113 78
rect 113 77 114 78
rect 6 76 7 77
rect 7 76 8 77
rect 8 76 9 77
rect 9 76 10 77
rect 10 76 11 77
rect 11 76 12 77
rect 12 76 13 77
rect 27 76 28 77
rect 28 76 29 77
rect 29 76 30 77
rect 30 76 31 77
rect 31 76 32 77
rect 32 76 33 77
rect 108 76 109 77
rect 109 76 110 77
rect 110 76 111 77
rect 111 76 112 77
rect 112 76 113 77
rect 113 76 114 77
rect 5 75 6 76
rect 6 75 7 76
rect 7 75 8 76
rect 8 75 9 76
rect 9 75 10 76
rect 27 75 28 76
rect 28 75 29 76
rect 29 75 30 76
rect 30 75 31 76
rect 31 75 32 76
rect 108 75 109 76
rect 109 75 110 76
rect 110 75 111 76
rect 111 75 112 76
rect 112 75 113 76
rect 113 75 114 76
rect 4 74 5 75
rect 5 74 6 75
rect 6 74 7 75
rect 7 74 8 75
rect 25 74 26 75
rect 26 74 27 75
rect 27 74 28 75
rect 28 74 29 75
rect 29 74 30 75
rect 30 74 31 75
rect 108 74 109 75
rect 109 74 110 75
rect 110 74 111 75
rect 111 74 112 75
rect 112 74 113 75
rect 113 74 114 75
rect 114 74 115 75
rect 4 73 5 74
rect 5 73 6 74
rect 6 73 7 74
rect 7 73 8 74
rect 25 73 26 74
rect 26 73 27 74
rect 27 73 28 74
rect 28 73 29 74
rect 29 73 30 74
rect 109 73 110 74
rect 110 73 111 74
rect 111 73 112 74
rect 112 73 113 74
rect 113 73 114 74
rect 114 73 115 74
rect 4 72 5 73
rect 5 72 6 73
rect 6 72 7 73
rect 7 72 8 73
rect 25 72 26 73
rect 26 72 27 73
rect 27 72 28 73
rect 28 72 29 73
rect 110 72 111 73
rect 111 72 112 73
rect 112 72 113 73
rect 113 72 114 73
rect 114 72 115 73
rect 4 71 5 72
rect 5 71 6 72
rect 6 71 7 72
rect 7 71 8 72
rect 24 71 25 72
rect 25 71 26 72
rect 26 71 27 72
rect 27 71 28 72
rect 110 71 111 72
rect 111 71 112 72
rect 112 71 113 72
rect 113 71 114 72
rect 114 71 115 72
rect 4 70 5 71
rect 5 70 6 71
rect 6 70 7 71
rect 7 70 8 71
rect 8 70 9 71
rect 23 70 24 71
rect 24 70 25 71
rect 25 70 26 71
rect 26 70 27 71
rect 27 70 28 71
rect 111 70 112 71
rect 112 70 113 71
rect 113 70 114 71
rect 114 70 115 71
rect 5 69 6 70
rect 6 69 7 70
rect 7 69 8 70
rect 8 69 9 70
rect 9 69 10 70
rect 23 69 24 70
rect 24 69 25 70
rect 25 69 26 70
rect 26 69 27 70
rect 111 69 112 70
rect 112 69 113 70
rect 113 69 114 70
rect 114 69 115 70
rect 5 68 6 69
rect 6 68 7 69
rect 7 68 8 69
rect 8 68 9 69
rect 9 68 10 69
rect 23 68 24 69
rect 24 68 25 69
rect 25 68 26 69
rect 112 68 113 69
rect 113 68 114 69
rect 114 68 115 69
rect 5 67 6 68
rect 6 67 7 68
rect 7 67 8 68
rect 8 67 9 68
rect 9 67 10 68
rect 10 67 11 68
rect 11 67 12 68
rect 22 67 23 68
rect 23 67 24 68
rect 24 67 25 68
rect 25 67 26 68
rect 112 67 113 68
rect 113 67 114 68
rect 114 67 115 68
rect 115 67 116 68
rect 7 66 8 67
rect 8 66 9 67
rect 9 66 10 67
rect 10 66 11 67
rect 11 66 12 67
rect 12 66 13 67
rect 22 66 23 67
rect 23 66 24 67
rect 24 66 25 67
rect 112 66 113 67
rect 113 66 114 67
rect 114 66 115 67
rect 115 66 116 67
rect 7 65 8 66
rect 8 65 9 66
rect 9 65 10 66
rect 10 65 11 66
rect 11 65 12 66
rect 12 65 13 66
rect 13 65 14 66
rect 21 65 22 66
rect 22 65 23 66
rect 23 65 24 66
rect 25 65 26 66
rect 26 65 27 66
rect 27 65 28 66
rect 28 65 29 66
rect 29 65 30 66
rect 30 65 31 66
rect 31 65 32 66
rect 32 65 33 66
rect 33 65 34 66
rect 34 65 35 66
rect 35 65 36 66
rect 36 65 37 66
rect 37 65 38 66
rect 112 65 113 66
rect 113 65 114 66
rect 114 65 115 66
rect 115 65 116 66
rect 9 64 10 65
rect 10 64 11 65
rect 11 64 12 65
rect 12 64 13 65
rect 13 64 14 65
rect 14 64 15 65
rect 15 64 16 65
rect 20 64 21 65
rect 21 64 22 65
rect 22 64 23 65
rect 23 64 24 65
rect 25 64 26 65
rect 26 64 27 65
rect 27 64 28 65
rect 28 64 29 65
rect 29 64 30 65
rect 30 64 31 65
rect 31 64 32 65
rect 32 64 33 65
rect 33 64 34 65
rect 34 64 35 65
rect 35 64 36 65
rect 36 64 37 65
rect 37 64 38 65
rect 113 64 114 65
rect 114 64 115 65
rect 115 64 116 65
rect 11 63 12 64
rect 12 63 13 64
rect 13 63 14 64
rect 14 63 15 64
rect 15 63 16 64
rect 16 63 17 64
rect 17 63 18 64
rect 18 63 19 64
rect 19 63 20 64
rect 20 63 21 64
rect 21 63 22 64
rect 22 63 23 64
rect 27 63 28 64
rect 28 63 29 64
rect 29 63 30 64
rect 33 63 34 64
rect 34 63 35 64
rect 35 63 36 64
rect 113 63 114 64
rect 114 63 115 64
rect 115 63 116 64
rect 13 62 14 63
rect 14 62 15 63
rect 15 62 16 63
rect 16 62 17 63
rect 17 62 18 63
rect 18 62 19 63
rect 19 62 20 63
rect 20 62 21 63
rect 21 62 22 63
rect 22 62 23 63
rect 27 62 28 63
rect 28 62 29 63
rect 29 62 30 63
rect 32 62 33 63
rect 33 62 34 63
rect 34 62 35 63
rect 113 62 114 63
rect 114 62 115 63
rect 115 62 116 63
rect 15 61 16 62
rect 16 61 17 62
rect 17 61 18 62
rect 18 61 19 62
rect 19 61 20 62
rect 20 61 21 62
rect 21 61 22 62
rect 27 61 28 62
rect 28 61 29 62
rect 29 61 30 62
rect 31 61 32 62
rect 32 61 33 62
rect 33 61 34 62
rect 113 61 114 62
rect 114 61 115 62
rect 115 61 116 62
rect 16 60 17 61
rect 17 60 18 61
rect 18 60 19 61
rect 19 60 20 61
rect 20 60 21 61
rect 21 60 22 61
rect 27 60 28 61
rect 28 60 29 61
rect 29 60 30 61
rect 30 60 31 61
rect 31 60 32 61
rect 32 60 33 61
rect 33 60 34 61
rect 100 60 101 61
rect 101 60 102 61
rect 102 60 103 61
rect 103 60 104 61
rect 104 60 105 61
rect 105 60 106 61
rect 106 60 107 61
rect 113 60 114 61
rect 114 60 115 61
rect 115 60 116 61
rect 18 59 19 60
rect 19 59 20 60
rect 20 59 21 60
rect 21 59 22 60
rect 27 59 28 60
rect 28 59 29 60
rect 29 59 30 60
rect 30 59 31 60
rect 31 59 32 60
rect 101 59 102 60
rect 102 59 103 60
rect 103 59 104 60
rect 104 59 105 60
rect 113 59 114 60
rect 114 59 115 60
rect 115 59 116 60
rect 19 58 20 59
rect 20 58 21 59
rect 21 58 22 59
rect 27 58 28 59
rect 28 58 29 59
rect 29 58 30 59
rect 30 58 31 59
rect 31 58 32 59
rect 32 58 33 59
rect 102 58 103 59
rect 103 58 104 59
rect 104 58 105 59
rect 113 58 114 59
rect 114 58 115 59
rect 115 58 116 59
rect 19 57 20 58
rect 20 57 21 58
rect 21 57 22 58
rect 27 57 28 58
rect 28 57 29 58
rect 29 57 30 58
rect 30 57 31 58
rect 31 57 32 58
rect 32 57 33 58
rect 33 57 34 58
rect 102 57 103 58
rect 103 57 104 58
rect 104 57 105 58
rect 113 57 114 58
rect 114 57 115 58
rect 115 57 116 58
rect 20 56 21 57
rect 27 56 28 57
rect 28 56 29 57
rect 29 56 30 57
rect 30 56 31 57
rect 31 56 32 57
rect 32 56 33 57
rect 33 56 34 57
rect 34 56 35 57
rect 41 56 42 57
rect 42 56 43 57
rect 102 56 103 57
rect 103 56 104 57
rect 104 56 105 57
rect 113 56 114 57
rect 114 56 115 57
rect 115 56 116 57
rect 20 55 21 56
rect 27 55 28 56
rect 28 55 29 56
rect 29 55 30 56
rect 31 55 32 56
rect 32 55 33 56
rect 33 55 34 56
rect 34 55 35 56
rect 35 55 36 56
rect 40 55 41 56
rect 41 55 42 56
rect 42 55 43 56
rect 102 55 103 56
rect 103 55 104 56
rect 104 55 105 56
rect 113 55 114 56
rect 114 55 115 56
rect 115 55 116 56
rect 20 54 21 55
rect 27 54 28 55
rect 28 54 29 55
rect 29 54 30 55
rect 32 54 33 55
rect 33 54 34 55
rect 34 54 35 55
rect 35 54 36 55
rect 40 54 41 55
rect 41 54 42 55
rect 42 54 43 55
rect 43 54 44 55
rect 102 54 103 55
rect 103 54 104 55
rect 104 54 105 55
rect 113 54 114 55
rect 114 54 115 55
rect 115 54 116 55
rect 20 53 21 54
rect 27 53 28 54
rect 28 53 29 54
rect 29 53 30 54
rect 33 53 34 54
rect 34 53 35 54
rect 35 53 36 54
rect 36 53 37 54
rect 39 53 40 54
rect 40 53 41 54
rect 41 53 42 54
rect 42 53 43 54
rect 43 53 44 54
rect 102 53 103 54
rect 103 53 104 54
rect 104 53 105 54
rect 113 53 114 54
rect 114 53 115 54
rect 115 53 116 54
rect 20 52 21 53
rect 27 52 28 53
rect 28 52 29 53
rect 29 52 30 53
rect 33 52 34 53
rect 34 52 35 53
rect 35 52 36 53
rect 36 52 37 53
rect 37 52 38 53
rect 39 52 40 53
rect 40 52 41 53
rect 41 52 42 53
rect 42 52 43 53
rect 43 52 44 53
rect 102 52 103 53
rect 103 52 104 53
rect 104 52 105 53
rect 113 52 114 53
rect 114 52 115 53
rect 19 51 20 52
rect 20 51 21 52
rect 25 51 26 52
rect 26 51 27 52
rect 27 51 28 52
rect 28 51 29 52
rect 29 51 30 52
rect 30 51 31 52
rect 32 51 33 52
rect 33 51 34 52
rect 34 51 35 52
rect 35 51 36 52
rect 36 51 37 52
rect 37 51 38 52
rect 38 51 39 52
rect 39 51 40 52
rect 40 51 41 52
rect 41 51 42 52
rect 42 51 43 52
rect 43 51 44 52
rect 44 51 45 52
rect 88 51 89 52
rect 89 51 90 52
rect 90 51 91 52
rect 91 51 92 52
rect 92 51 93 52
rect 93 51 94 52
rect 94 51 95 52
rect 95 51 96 52
rect 96 51 97 52
rect 97 51 98 52
rect 98 51 99 52
rect 99 51 100 52
rect 102 51 103 52
rect 103 51 104 52
rect 104 51 105 52
rect 112 51 113 52
rect 113 51 114 52
rect 114 51 115 52
rect 19 50 20 51
rect 20 50 21 51
rect 38 50 39 51
rect 39 50 40 51
rect 41 50 42 51
rect 42 50 43 51
rect 43 50 44 51
rect 44 50 45 51
rect 88 50 89 51
rect 89 50 90 51
rect 90 50 91 51
rect 91 50 92 51
rect 92 50 93 51
rect 93 50 94 51
rect 94 50 95 51
rect 95 50 96 51
rect 96 50 97 51
rect 97 50 98 51
rect 98 50 99 51
rect 99 50 100 51
rect 100 50 101 51
rect 102 50 103 51
rect 103 50 104 51
rect 104 50 105 51
rect 112 50 113 51
rect 113 50 114 51
rect 114 50 115 51
rect 19 49 20 50
rect 20 49 21 50
rect 21 49 22 50
rect 38 49 39 50
rect 39 49 40 50
rect 42 49 43 50
rect 43 49 44 50
rect 44 49 45 50
rect 88 49 89 50
rect 89 49 90 50
rect 90 49 91 50
rect 91 49 92 50
rect 92 49 93 50
rect 93 49 94 50
rect 94 49 95 50
rect 95 49 96 50
rect 96 49 97 50
rect 97 49 98 50
rect 98 49 99 50
rect 99 49 100 50
rect 102 49 103 50
rect 103 49 104 50
rect 104 49 105 50
rect 112 49 113 50
rect 113 49 114 50
rect 114 49 115 50
rect 19 48 20 49
rect 20 48 21 49
rect 21 48 22 49
rect 37 48 38 49
rect 38 48 39 49
rect 39 48 40 49
rect 40 48 41 49
rect 41 48 42 49
rect 42 48 43 49
rect 43 48 44 49
rect 44 48 45 49
rect 45 48 46 49
rect 88 48 89 49
rect 89 48 90 49
rect 90 48 91 49
rect 92 48 93 49
rect 93 48 94 49
rect 94 48 95 49
rect 95 48 96 49
rect 98 48 99 49
rect 99 48 100 49
rect 100 48 101 49
rect 102 48 103 49
rect 103 48 104 49
rect 104 48 105 49
rect 112 48 113 49
rect 113 48 114 49
rect 114 48 115 49
rect 19 47 20 48
rect 20 47 21 48
rect 21 47 22 48
rect 37 47 38 48
rect 38 47 39 48
rect 39 47 40 48
rect 40 47 41 48
rect 41 47 42 48
rect 42 47 43 48
rect 43 47 44 48
rect 44 47 45 48
rect 45 47 46 48
rect 88 47 89 48
rect 89 47 90 48
rect 93 47 94 48
rect 94 47 95 48
rect 95 47 96 48
rect 98 47 99 48
rect 99 47 100 48
rect 100 47 101 48
rect 101 47 102 48
rect 102 47 103 48
rect 103 47 104 48
rect 104 47 105 48
rect 105 47 106 48
rect 106 47 107 48
rect 112 47 113 48
rect 113 47 114 48
rect 114 47 115 48
rect 19 46 20 47
rect 20 46 21 47
rect 21 46 22 47
rect 37 46 38 47
rect 38 46 39 47
rect 43 46 44 47
rect 44 46 45 47
rect 45 46 46 47
rect 92 46 93 47
rect 93 46 94 47
rect 94 46 95 47
rect 95 46 96 47
rect 100 46 101 47
rect 101 46 102 47
rect 102 46 103 47
rect 103 46 104 47
rect 104 46 105 47
rect 105 46 106 47
rect 106 46 107 47
rect 111 46 112 47
rect 112 46 113 47
rect 113 46 114 47
rect 114 46 115 47
rect 19 45 20 46
rect 20 45 21 46
rect 21 45 22 46
rect 36 45 37 46
rect 37 45 38 46
rect 38 45 39 46
rect 43 45 44 46
rect 44 45 45 46
rect 45 45 46 46
rect 46 45 47 46
rect 92 45 93 46
rect 93 45 94 46
rect 94 45 95 46
rect 95 45 96 46
rect 111 45 112 46
rect 112 45 113 46
rect 113 45 114 46
rect 19 44 20 45
rect 20 44 21 45
rect 21 44 22 45
rect 36 44 37 45
rect 37 44 38 45
rect 44 44 45 45
rect 45 44 46 45
rect 46 44 47 45
rect 48 44 49 45
rect 49 44 50 45
rect 92 44 93 45
rect 93 44 94 45
rect 94 44 95 45
rect 95 44 96 45
rect 110 44 111 45
rect 111 44 112 45
rect 112 44 113 45
rect 113 44 114 45
rect 20 43 21 44
rect 21 43 22 44
rect 22 43 23 44
rect 35 43 36 44
rect 36 43 37 44
rect 37 43 38 44
rect 38 43 39 44
rect 43 43 44 44
rect 44 43 45 44
rect 45 43 46 44
rect 46 43 47 44
rect 47 43 48 44
rect 48 43 49 44
rect 49 43 50 44
rect 77 43 78 44
rect 78 43 79 44
rect 79 43 80 44
rect 80 43 81 44
rect 81 43 82 44
rect 82 43 83 44
rect 83 43 84 44
rect 84 43 85 44
rect 85 43 86 44
rect 86 43 87 44
rect 87 43 88 44
rect 92 43 93 44
rect 93 43 94 44
rect 94 43 95 44
rect 95 43 96 44
rect 110 43 111 44
rect 111 43 112 44
rect 112 43 113 44
rect 113 43 114 44
rect 20 42 21 43
rect 21 42 22 43
rect 22 42 23 43
rect 35 42 36 43
rect 36 42 37 43
rect 37 42 38 43
rect 38 42 39 43
rect 43 42 44 43
rect 44 42 45 43
rect 45 42 46 43
rect 46 42 47 43
rect 47 42 48 43
rect 48 42 49 43
rect 49 42 50 43
rect 77 42 78 43
rect 78 42 79 43
rect 79 42 80 43
rect 80 42 81 43
rect 81 42 82 43
rect 82 42 83 43
rect 83 42 84 43
rect 84 42 85 43
rect 85 42 86 43
rect 86 42 87 43
rect 87 42 88 43
rect 92 42 93 43
rect 93 42 94 43
rect 94 42 95 43
rect 95 42 96 43
rect 110 42 111 43
rect 111 42 112 43
rect 112 42 113 43
rect 20 41 21 42
rect 21 41 22 42
rect 22 41 23 42
rect 47 41 48 42
rect 48 41 49 42
rect 49 41 50 42
rect 50 41 51 42
rect 62 41 63 42
rect 77 41 78 42
rect 78 41 79 42
rect 79 41 80 42
rect 80 41 81 42
rect 81 41 82 42
rect 82 41 83 42
rect 83 41 84 42
rect 84 41 85 42
rect 85 41 86 42
rect 86 41 87 42
rect 87 41 88 42
rect 92 41 93 42
rect 93 41 94 42
rect 94 41 95 42
rect 95 41 96 42
rect 109 41 110 42
rect 110 41 111 42
rect 111 41 112 42
rect 112 41 113 42
rect 21 40 22 41
rect 22 40 23 41
rect 23 40 24 41
rect 47 40 48 41
rect 48 40 49 41
rect 49 40 50 41
rect 50 40 51 41
rect 61 40 62 41
rect 62 40 63 41
rect 63 40 64 41
rect 78 40 79 41
rect 79 40 80 41
rect 80 40 81 41
rect 81 40 82 41
rect 82 40 83 41
rect 86 40 87 41
rect 87 40 88 41
rect 92 40 93 41
rect 93 40 94 41
rect 94 40 95 41
rect 95 40 96 41
rect 108 40 109 41
rect 109 40 110 41
rect 110 40 111 41
rect 111 40 112 41
rect 112 40 113 41
rect 21 39 22 40
rect 22 39 23 40
rect 23 39 24 40
rect 46 39 47 40
rect 47 39 48 40
rect 48 39 49 40
rect 49 39 50 40
rect 50 39 51 40
rect 51 39 52 40
rect 61 39 62 40
rect 62 39 63 40
rect 63 39 64 40
rect 79 39 80 40
rect 80 39 81 40
rect 81 39 82 40
rect 82 39 83 40
rect 86 39 87 40
rect 87 39 88 40
rect 92 39 93 40
rect 93 39 94 40
rect 94 39 95 40
rect 95 39 96 40
rect 108 39 109 40
rect 109 39 110 40
rect 110 39 111 40
rect 111 39 112 40
rect 112 39 113 40
rect 21 38 22 39
rect 22 38 23 39
rect 23 38 24 39
rect 46 38 47 39
rect 47 38 48 39
rect 48 38 49 39
rect 49 38 50 39
rect 50 38 51 39
rect 51 38 52 39
rect 61 38 62 39
rect 62 38 63 39
rect 63 38 64 39
rect 64 38 65 39
rect 70 38 71 39
rect 71 38 72 39
rect 72 38 73 39
rect 73 38 74 39
rect 74 38 75 39
rect 75 38 76 39
rect 79 38 80 39
rect 80 38 81 39
rect 81 38 82 39
rect 82 38 83 39
rect 83 38 84 39
rect 92 38 93 39
rect 93 38 94 39
rect 94 38 95 39
rect 95 38 96 39
rect 108 38 109 39
rect 109 38 110 39
rect 110 38 111 39
rect 111 38 112 39
rect 21 37 22 38
rect 22 37 23 38
rect 23 37 24 38
rect 24 37 25 38
rect 45 37 46 38
rect 46 37 47 38
rect 47 37 48 38
rect 49 37 50 38
rect 50 37 51 38
rect 51 37 52 38
rect 60 37 61 38
rect 61 37 62 38
rect 62 37 63 38
rect 63 37 64 38
rect 64 37 65 38
rect 71 37 72 38
rect 72 37 73 38
rect 73 37 74 38
rect 74 37 75 38
rect 75 37 76 38
rect 80 37 81 38
rect 81 37 82 38
rect 82 37 83 38
rect 83 37 84 38
rect 84 37 85 38
rect 91 37 92 38
rect 92 37 93 38
rect 93 37 94 38
rect 94 37 95 38
rect 95 37 96 38
rect 96 37 97 38
rect 97 37 98 38
rect 107 37 108 38
rect 108 37 109 38
rect 109 37 110 38
rect 110 37 111 38
rect 111 37 112 38
rect 22 36 23 37
rect 23 36 24 37
rect 24 36 25 37
rect 45 36 46 37
rect 46 36 47 37
rect 49 36 50 37
rect 50 36 51 37
rect 51 36 52 37
rect 52 36 53 37
rect 60 36 61 37
rect 61 36 62 37
rect 62 36 63 37
rect 63 36 64 37
rect 64 36 65 37
rect 72 36 73 37
rect 73 36 74 37
rect 74 36 75 37
rect 81 36 82 37
rect 82 36 83 37
rect 83 36 84 37
rect 84 36 85 37
rect 91 36 92 37
rect 92 36 93 37
rect 93 36 94 37
rect 94 36 95 37
rect 95 36 96 37
rect 96 36 97 37
rect 97 36 98 37
rect 106 36 107 37
rect 107 36 108 37
rect 108 36 109 37
rect 109 36 110 37
rect 110 36 111 37
rect 22 35 23 36
rect 23 35 24 36
rect 24 35 25 36
rect 25 35 26 36
rect 45 35 46 36
rect 46 35 47 36
rect 49 35 50 36
rect 50 35 51 36
rect 51 35 52 36
rect 52 35 53 36
rect 59 35 60 36
rect 60 35 61 36
rect 61 35 62 36
rect 62 35 63 36
rect 63 35 64 36
rect 64 35 65 36
rect 65 35 66 36
rect 72 35 73 36
rect 73 35 74 36
rect 74 35 75 36
rect 81 35 82 36
rect 82 35 83 36
rect 83 35 84 36
rect 106 35 107 36
rect 107 35 108 36
rect 108 35 109 36
rect 109 35 110 36
rect 110 35 111 36
rect 23 34 24 35
rect 24 34 25 35
rect 25 34 26 35
rect 44 34 45 35
rect 45 34 46 35
rect 46 34 47 35
rect 50 34 51 35
rect 51 34 52 35
rect 52 34 53 35
rect 53 34 54 35
rect 59 34 60 35
rect 60 34 61 35
rect 61 34 62 35
rect 62 34 63 35
rect 63 34 64 35
rect 64 34 65 35
rect 65 34 66 35
rect 72 34 73 35
rect 73 34 74 35
rect 74 34 75 35
rect 80 34 81 35
rect 81 34 82 35
rect 82 34 83 35
rect 83 34 84 35
rect 104 34 105 35
rect 105 34 106 35
rect 106 34 107 35
rect 107 34 108 35
rect 108 34 109 35
rect 109 34 110 35
rect 110 34 111 35
rect 23 33 24 34
rect 24 33 25 34
rect 25 33 26 34
rect 44 33 45 34
rect 45 33 46 34
rect 50 33 51 34
rect 51 33 52 34
rect 52 33 53 34
rect 53 33 54 34
rect 59 33 60 34
rect 60 33 61 34
rect 63 33 64 34
rect 64 33 65 34
rect 65 33 66 34
rect 66 33 67 34
rect 72 33 73 34
rect 73 33 74 34
rect 74 33 75 34
rect 80 33 81 34
rect 81 33 82 34
rect 82 33 83 34
rect 87 33 88 34
rect 88 33 89 34
rect 104 33 105 34
rect 105 33 106 34
rect 106 33 107 34
rect 107 33 108 34
rect 108 33 109 34
rect 109 33 110 34
rect 23 32 24 33
rect 24 32 25 33
rect 25 32 26 33
rect 26 32 27 33
rect 44 32 45 33
rect 45 32 46 33
rect 51 32 52 33
rect 52 32 53 33
rect 53 32 54 33
rect 58 32 59 33
rect 59 32 60 33
rect 60 32 61 33
rect 63 32 64 33
rect 64 32 65 33
rect 65 32 66 33
rect 66 32 67 33
rect 72 32 73 33
rect 73 32 74 33
rect 74 32 75 33
rect 79 32 80 33
rect 80 32 81 33
rect 81 32 82 33
rect 87 32 88 33
rect 88 32 89 33
rect 103 32 104 33
rect 104 32 105 33
rect 105 32 106 33
rect 106 32 107 33
rect 107 32 108 33
rect 108 32 109 33
rect 24 31 25 32
rect 25 31 26 32
rect 26 31 27 32
rect 27 31 28 32
rect 42 31 43 32
rect 43 31 44 32
rect 44 31 45 32
rect 45 31 46 32
rect 46 31 47 32
rect 49 31 50 32
rect 50 31 51 32
rect 51 31 52 32
rect 52 31 53 32
rect 53 31 54 32
rect 54 31 55 32
rect 55 31 56 32
rect 58 31 59 32
rect 59 31 60 32
rect 64 31 65 32
rect 65 31 66 32
rect 66 31 67 32
rect 72 31 73 32
rect 73 31 74 32
rect 74 31 75 32
rect 78 31 79 32
rect 79 31 80 32
rect 80 31 81 32
rect 81 31 82 32
rect 82 31 83 32
rect 83 31 84 32
rect 84 31 85 32
rect 85 31 86 32
rect 86 31 87 32
rect 87 31 88 32
rect 88 31 89 32
rect 102 31 103 32
rect 103 31 104 32
rect 104 31 105 32
rect 105 31 106 32
rect 106 31 107 32
rect 107 31 108 32
rect 24 30 25 31
rect 25 30 26 31
rect 26 30 27 31
rect 27 30 28 31
rect 42 30 43 31
rect 43 30 44 31
rect 44 30 45 31
rect 45 30 46 31
rect 46 30 47 31
rect 49 30 50 31
rect 50 30 51 31
rect 51 30 52 31
rect 52 30 53 31
rect 53 30 54 31
rect 54 30 55 31
rect 55 30 56 31
rect 58 30 59 31
rect 59 30 60 31
rect 64 30 65 31
rect 65 30 66 31
rect 66 30 67 31
rect 67 30 68 31
rect 72 30 73 31
rect 73 30 74 31
rect 74 30 75 31
rect 77 30 78 31
rect 78 30 79 31
rect 79 30 80 31
rect 80 30 81 31
rect 81 30 82 31
rect 82 30 83 31
rect 83 30 84 31
rect 84 30 85 31
rect 85 30 86 31
rect 86 30 87 31
rect 87 30 88 31
rect 101 30 102 31
rect 102 30 103 31
rect 103 30 104 31
rect 104 30 105 31
rect 105 30 106 31
rect 106 30 107 31
rect 25 29 26 30
rect 26 29 27 30
rect 27 29 28 30
rect 28 29 29 30
rect 57 29 58 30
rect 58 29 59 30
rect 59 29 60 30
rect 64 29 65 30
rect 65 29 66 30
rect 66 29 67 30
rect 67 29 68 30
rect 72 29 73 30
rect 73 29 74 30
rect 74 29 75 30
rect 76 29 77 30
rect 77 29 78 30
rect 78 29 79 30
rect 79 29 80 30
rect 80 29 81 30
rect 81 29 82 30
rect 82 29 83 30
rect 83 29 84 30
rect 84 29 85 30
rect 85 29 86 30
rect 86 29 87 30
rect 87 29 88 30
rect 100 29 101 30
rect 101 29 102 30
rect 102 29 103 30
rect 103 29 104 30
rect 104 29 105 30
rect 105 29 106 30
rect 106 29 107 30
rect 25 28 26 29
rect 26 28 27 29
rect 27 28 28 29
rect 28 28 29 29
rect 56 28 57 29
rect 57 28 58 29
rect 58 28 59 29
rect 59 28 60 29
rect 64 28 65 29
rect 65 28 66 29
rect 66 28 67 29
rect 67 28 68 29
rect 68 28 69 29
rect 72 28 73 29
rect 73 28 74 29
rect 74 28 75 29
rect 76 28 77 29
rect 77 28 78 29
rect 78 28 79 29
rect 79 28 80 29
rect 80 28 81 29
rect 81 28 82 29
rect 82 28 83 29
rect 83 28 84 29
rect 84 28 85 29
rect 85 28 86 29
rect 86 28 87 29
rect 87 28 88 29
rect 99 28 100 29
rect 100 28 101 29
rect 101 28 102 29
rect 102 28 103 29
rect 103 28 104 29
rect 104 28 105 29
rect 105 28 106 29
rect 26 27 27 28
rect 27 27 28 28
rect 28 27 29 28
rect 29 27 30 28
rect 55 27 56 28
rect 56 27 57 28
rect 57 27 58 28
rect 58 27 59 28
rect 59 27 60 28
rect 60 27 61 28
rect 63 27 64 28
rect 64 27 65 28
rect 65 27 66 28
rect 66 27 67 28
rect 67 27 68 28
rect 68 27 69 28
rect 69 27 70 28
rect 72 27 73 28
rect 73 27 74 28
rect 74 27 75 28
rect 98 27 99 28
rect 99 27 100 28
rect 100 27 101 28
rect 101 27 102 28
rect 102 27 103 28
rect 103 27 104 28
rect 104 27 105 28
rect 27 26 28 27
rect 28 26 29 27
rect 29 26 30 27
rect 30 26 31 27
rect 72 26 73 27
rect 73 26 74 27
rect 74 26 75 27
rect 97 26 98 27
rect 98 26 99 27
rect 99 26 100 27
rect 100 26 101 27
rect 101 26 102 27
rect 102 26 103 27
rect 27 25 28 26
rect 28 25 29 26
rect 29 25 30 26
rect 30 25 31 26
rect 31 25 32 26
rect 71 25 72 26
rect 72 25 73 26
rect 73 25 74 26
rect 74 25 75 26
rect 96 25 97 26
rect 97 25 98 26
rect 98 25 99 26
rect 99 25 100 26
rect 100 25 101 26
rect 101 25 102 26
rect 102 25 103 26
rect 28 24 29 25
rect 29 24 30 25
rect 30 24 31 25
rect 31 24 32 25
rect 70 24 71 25
rect 71 24 72 25
rect 72 24 73 25
rect 73 24 74 25
rect 74 24 75 25
rect 75 24 76 25
rect 94 24 95 25
rect 95 24 96 25
rect 96 24 97 25
rect 97 24 98 25
rect 98 24 99 25
rect 99 24 100 25
rect 100 24 101 25
rect 101 24 102 25
rect 29 23 30 24
rect 30 23 31 24
rect 31 23 32 24
rect 32 23 33 24
rect 93 23 94 24
rect 94 23 95 24
rect 95 23 96 24
rect 96 23 97 24
rect 97 23 98 24
rect 98 23 99 24
rect 99 23 100 24
rect 29 22 30 23
rect 30 22 31 23
rect 31 22 32 23
rect 32 22 33 23
rect 33 22 34 23
rect 92 22 93 23
rect 93 22 94 23
rect 94 22 95 23
rect 95 22 96 23
rect 96 22 97 23
rect 97 22 98 23
rect 98 22 99 23
rect 30 21 31 22
rect 31 21 32 22
rect 32 21 33 22
rect 33 21 34 22
rect 34 21 35 22
rect 91 21 92 22
rect 92 21 93 22
rect 93 21 94 22
rect 94 21 95 22
rect 95 21 96 22
rect 96 21 97 22
rect 97 21 98 22
rect 31 20 32 21
rect 32 20 33 21
rect 33 20 34 21
rect 34 20 35 21
rect 35 20 36 21
rect 90 20 91 21
rect 91 20 92 21
rect 92 20 93 21
rect 93 20 94 21
rect 94 20 95 21
rect 95 20 96 21
rect 96 20 97 21
rect 32 19 33 20
rect 33 19 34 20
rect 34 19 35 20
rect 35 19 36 20
rect 36 19 37 20
rect 90 19 91 20
rect 91 19 92 20
rect 92 19 93 20
rect 93 19 94 20
rect 94 19 95 20
rect 33 18 34 19
rect 34 18 35 19
rect 35 18 36 19
rect 36 18 37 19
rect 37 18 38 19
rect 38 18 39 19
rect 88 18 89 19
rect 89 18 90 19
rect 90 18 91 19
rect 91 18 92 19
rect 92 18 93 19
rect 93 18 94 19
rect 94 18 95 19
rect 34 17 35 18
rect 35 17 36 18
rect 36 17 37 18
rect 37 17 38 18
rect 38 17 39 18
rect 39 17 40 18
rect 87 17 88 18
rect 88 17 89 18
rect 89 17 90 18
rect 90 17 91 18
rect 91 17 92 18
rect 92 17 93 18
rect 35 16 36 17
rect 36 16 37 17
rect 37 16 38 17
rect 38 16 39 17
rect 39 16 40 17
rect 40 16 41 17
rect 86 16 87 17
rect 87 16 88 17
rect 88 16 89 17
rect 89 16 90 17
rect 90 16 91 17
rect 36 15 37 16
rect 37 15 38 16
rect 38 15 39 16
rect 39 15 40 16
rect 40 15 41 16
rect 41 15 42 16
rect 86 15 87 16
rect 87 15 88 16
rect 88 15 89 16
rect 89 15 90 16
rect 37 14 38 15
rect 38 14 39 15
rect 39 14 40 15
rect 40 14 41 15
rect 41 14 42 15
rect 42 14 43 15
rect 43 14 44 15
rect 68 14 69 15
rect 69 14 70 15
rect 84 14 85 15
rect 85 14 86 15
rect 86 14 87 15
rect 87 14 88 15
rect 88 14 89 15
rect 39 13 40 14
rect 40 13 41 14
rect 41 13 42 14
rect 42 13 43 14
rect 43 13 44 14
rect 44 13 45 14
rect 45 13 46 14
rect 46 13 47 14
rect 47 13 48 14
rect 48 13 49 14
rect 64 13 65 14
rect 65 13 66 14
rect 66 13 67 14
rect 67 13 68 14
rect 68 13 69 14
rect 69 13 70 14
rect 83 13 84 14
rect 84 13 85 14
rect 85 13 86 14
rect 86 13 87 14
rect 40 12 41 13
rect 41 12 42 13
rect 42 12 43 13
rect 43 12 44 13
rect 44 12 45 13
rect 45 12 46 13
rect 46 12 47 13
rect 47 12 48 13
rect 48 12 49 13
rect 49 12 50 13
rect 50 12 51 13
rect 51 12 52 13
rect 52 12 53 13
rect 53 12 54 13
rect 54 12 55 13
rect 55 12 56 13
rect 56 12 57 13
rect 57 12 58 13
rect 58 12 59 13
rect 59 12 60 13
rect 60 12 61 13
rect 61 12 62 13
rect 62 12 63 13
rect 63 12 64 13
rect 64 12 65 13
rect 65 12 66 13
rect 66 12 67 13
rect 67 12 68 13
rect 68 12 69 13
rect 82 12 83 13
rect 83 12 84 13
rect 84 12 85 13
rect 85 12 86 13
rect 41 11 42 12
rect 42 11 43 12
rect 43 11 44 12
rect 44 11 45 12
rect 45 11 46 12
rect 46 11 47 12
rect 47 11 48 12
rect 48 11 49 12
rect 49 11 50 12
rect 50 11 51 12
rect 51 11 52 12
rect 52 11 53 12
rect 53 11 54 12
rect 54 11 55 12
rect 55 11 56 12
rect 56 11 57 12
rect 57 11 58 12
rect 58 11 59 12
rect 59 11 60 12
rect 60 11 61 12
rect 61 11 62 12
rect 62 11 63 12
rect 63 11 64 12
rect 64 11 65 12
rect 65 11 66 12
rect 66 11 67 12
rect 67 11 68 12
rect 80 11 81 12
rect 81 11 82 12
rect 82 11 83 12
rect 83 11 84 12
rect 84 11 85 12
rect 44 10 45 11
rect 45 10 46 11
rect 46 10 47 11
rect 47 10 48 11
rect 48 10 49 11
rect 49 10 50 11
rect 50 10 51 11
rect 51 10 52 11
rect 52 10 53 11
rect 53 10 54 11
rect 54 10 55 11
rect 55 10 56 11
rect 56 10 57 11
rect 57 10 58 11
rect 58 10 59 11
rect 59 10 60 11
rect 60 10 61 11
rect 61 10 62 11
rect 62 10 63 11
rect 63 10 64 11
rect 64 10 65 11
rect 65 10 66 11
rect 66 10 67 11
rect 67 10 68 11
rect 68 10 69 11
rect 69 10 70 11
rect 78 10 79 11
rect 79 10 80 11
rect 80 10 81 11
rect 81 10 82 11
rect 82 10 83 11
rect 45 9 46 10
rect 46 9 47 10
rect 54 9 55 10
rect 55 9 56 10
rect 56 9 57 10
rect 57 9 58 10
rect 58 9 59 10
rect 59 9 60 10
rect 60 9 61 10
rect 61 9 62 10
rect 62 9 63 10
rect 63 9 64 10
rect 64 9 65 10
rect 65 9 66 10
rect 66 9 67 10
rect 67 9 68 10
rect 68 9 69 10
rect 69 9 70 10
rect 70 9 71 10
rect 71 9 72 10
rect 72 9 73 10
rect 73 9 74 10
rect 74 9 75 10
rect 75 9 76 10
rect 76 9 77 10
rect 77 9 78 10
rect 78 9 79 10
rect 79 9 80 10
rect 80 9 81 10
rect 81 9 82 10
rect 57 8 58 9
rect 58 8 59 9
rect 59 8 60 9
rect 60 8 61 9
rect 61 8 62 9
rect 62 8 63 9
rect 63 8 64 9
rect 64 8 65 9
rect 65 8 66 9
rect 66 8 67 9
rect 67 8 68 9
rect 68 8 69 9
rect 69 8 70 9
rect 70 8 71 9
rect 71 8 72 9
rect 72 8 73 9
rect 73 8 74 9
rect 74 8 75 9
rect 75 8 76 9
rect 76 8 77 9
rect 77 8 78 9
rect 78 8 79 9
rect 79 8 80 9
rect 80 8 81 9
rect 61 7 62 8
rect 62 7 63 8
rect 63 7 64 8
rect 64 7 65 8
rect 65 7 66 8
rect 66 7 67 8
rect 67 7 68 8
rect 68 7 69 8
rect 69 7 70 8
rect 70 7 71 8
rect 71 7 72 8
rect 72 7 73 8
rect 73 7 74 8
rect 74 7 75 8
rect 75 7 76 8
rect 76 7 77 8
rect 77 7 78 8
rect 78 7 79 8
rect 64 6 65 7
rect 65 6 66 7
rect 66 6 67 7
rect 67 6 68 7
rect 68 6 69 7
rect 69 6 70 7
rect 70 6 71 7
rect 71 6 72 7
rect 72 6 73 7
rect 73 6 74 7
rect 74 6 75 7
rect 75 6 76 7
rect 76 6 77 7
rect 77 6 78 7
rect 66 5 67 6
rect 67 5 68 6
rect 68 5 69 6
rect 69 5 70 6
rect 70 5 71 6
rect 71 5 72 6
rect 72 5 73 6
rect 73 5 74 6
rect 74 5 75 6
rect 75 5 76 6
rect 76 5 77 6
rect 70 4 71 5
rect 71 4 72 5
rect 72 4 73 5
rect 73 4 74 5
rect 74 4 75 5
rect 75 4 76 5
<< end >>
