magic
tech scmos
timestamp 1539608411
<< nwell >>
rect 116 172 184 184
rect 116 128 128 172
rect 172 128 184 172
rect 116 116 184 128
<< metal1 >>
rect 100 208 200 218
rect 145 182 155 208
rect 118 180 182 182
rect 118 176 120 180
rect 124 176 128 180
rect 132 176 136 180
rect 140 176 144 180
rect 148 176 152 180
rect 156 176 160 180
rect 164 176 168 180
rect 172 176 176 180
rect 180 176 182 180
rect 118 174 182 176
rect 118 172 126 174
rect 118 168 120 172
rect 124 168 126 172
rect 174 172 182 174
rect 118 164 126 168
rect 118 160 120 164
rect 124 160 126 164
rect 118 156 126 160
rect 118 152 120 156
rect 124 152 126 156
rect 118 148 126 152
rect 118 144 120 148
rect 124 144 126 148
rect 118 140 126 144
rect 118 136 120 140
rect 124 136 126 140
rect 118 132 126 136
rect 118 128 120 132
rect 124 128 126 132
rect 130 162 170 170
rect 130 130 138 162
rect 142 142 158 158
rect 118 124 126 128
rect 118 120 120 124
rect 124 120 126 124
rect 118 118 126 120
rect 142 85 152 142
rect 100 75 152 85
rect 162 90 170 162
rect 174 168 176 172
rect 180 168 182 172
rect 174 164 182 168
rect 174 160 176 164
rect 180 160 182 164
rect 174 156 182 160
rect 174 152 176 156
rect 180 152 182 156
rect 174 148 182 152
rect 174 144 176 148
rect 180 144 182 148
rect 174 140 182 144
rect 174 136 176 140
rect 180 136 182 140
rect 174 132 182 136
rect 174 128 176 132
rect 180 128 182 132
rect 174 124 182 128
rect 174 120 176 124
rect 180 120 182 124
rect 174 118 182 120
rect 162 80 200 90
<< pbase >>
rect 128 160 172 172
rect 128 140 140 160
rect 160 140 172 160
rect 128 128 172 140
<< nwpnbase >>
rect 140 140 160 160
<< pbasepdiffcontact >>
rect 132 164 136 168
rect 140 164 144 168
rect 156 164 160 168
rect 164 164 168 168
rect 132 156 136 160
rect 164 156 168 160
rect 132 140 136 144
rect 164 140 168 144
rect 132 132 136 136
rect 164 132 168 136
<< nbasendiffcontact >>
rect 144 152 148 156
rect 152 152 156 156
rect 144 144 148 148
rect 152 144 156 148
<< pdcontact >>
rect 120 176 124 180
rect 128 176 132 180
rect 136 176 140 180
rect 144 176 148 180
rect 152 176 156 180
rect 160 176 164 180
rect 168 176 172 180
rect 176 176 180 180
rect 120 168 124 172
rect 176 168 180 172
rect 120 160 124 164
rect 176 160 180 164
rect 120 152 124 156
rect 176 152 180 156
rect 120 144 124 148
rect 176 144 180 148
rect 120 136 124 140
rect 176 136 180 140
rect 120 128 124 132
rect 176 128 180 132
rect 120 120 124 124
rect 176 120 180 124
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_CHAR_c  L500_CHAR_c_0
timestamp 1534321654
transform 1 0 146 0 1 218
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_CHAR_n  L500_CHAR_n_0
timestamp 1534323117
transform 1 0 208 0 1 136
box 0 0 12 18
use L500_CHAR_p  L500_CHAR_p_0
timestamp 1534323210
transform 1 0 221 0 1 136
box 0 0 12 18
use L500_CHAR_n  L500_CHAR_n_0
timestamp 1534323117
transform 1 0 234 0 1 136
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_CHAR_e  L500_CHAR_e_0
timestamp 1534321786
transform 1 0 114 0 1 57
box 0 0 12 18
use L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 173 0 1 63
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
