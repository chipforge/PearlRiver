magic
tech scmos
timestamp 1540534746
<< polysilicon >>
rect 140 176 160 199
rect 140 102 160 125
<< metal1 >>
rect 100 225 200 245
rect 140 219 160 225
rect 140 75 160 82
rect 100 55 200 75
<< rndiffusion >>
rect 140 153 160 176
<< rpdiffusion >>
rect 140 125 160 148
<< rpoly >>
rect 140 148 160 153
<< polycontact >>
rect 140 199 160 219
rect 140 82 160 102
use L500_TPAD_blank  L500_TPAD_blank_2 ./Library/magic
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
