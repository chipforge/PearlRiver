magic
tech scmos
timestamp 1539768844
<< polysilicon >>
rect 145 165 155 171
rect 145 129 155 135
<< metal1 >>
rect 90 181 100 200
rect 200 181 210 200
rect 90 171 145 181
rect 155 171 210 181
rect 90 119 145 129
rect 155 119 210 129
rect 90 100 100 119
rect 200 100 210 119
<< rndiffusion >>
rect 145 153 155 159
<< rpdiffusion >>
rect 145 141 155 147
<< rpoly >>
rect 145 147 155 153
<< polycontact >>
rect 145 171 155 181
rect 145 119 155 129
<< polyndiff >>
rect 145 159 155 165
<< polypdiff >>
rect 145 135 155 141
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
