magic
tech scmos
timestamp 1541105161
<< error_s >>
rect 179 174 193 179
rect 130 170 131 171
rect 169 170 170 171
rect 129 169 171 170
rect 130 166 170 169
rect 130 134 134 166
rect 140 156 160 160
rect 140 144 144 156
rect 156 144 160 156
rect 140 140 160 144
rect 166 134 170 166
rect 130 130 170 134
rect 184 127 185 174
rect 188 127 193 174
rect 184 126 193 127
rect 122 122 178 124
rect 112 112 188 114
<< nwell >>
rect 106 178 194 194
rect 106 122 122 178
rect 134 160 166 166
rect 134 140 140 160
rect 160 140 166 160
rect 134 134 166 140
rect 178 122 194 178
rect 106 114 194 122
<< metal1 >>
rect 100 208 200 218
rect 145 176 155 208
rect 124 174 176 176
rect 124 126 126 174
rect 130 168 170 170
rect 130 126 132 168
rect 124 124 132 126
rect 142 142 158 158
rect 142 85 152 142
rect 168 126 170 168
rect 174 126 176 174
rect 168 124 176 126
rect 182 174 190 176
rect 182 126 184 174
rect 188 126 190 174
rect 100 75 152 85
rect 182 90 190 126
rect 182 80 200 90
<< nwpbase >>
rect 122 166 178 178
rect 122 134 134 166
rect 140 140 160 160
rect 166 134 178 166
rect 122 122 178 134
<< pbasepdiffcontact >>
rect 144 152 148 156
rect 152 152 156 156
rect 144 144 148 148
rect 152 144 156 148
<< ndcontact >>
rect 184 126 188 174
<< pdcontact >>
rect 126 170 174 174
rect 126 126 130 170
rect 170 126 174 170
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_CHAR_c  L500_CHAR_c_0
timestamp 1534321654
transform 1 0 146 0 1 230
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_CHAR_p  L500_CHAR_p_0
timestamp 1534323210
transform 1 0 208 0 1 136
box 0 0 12 18
use L500_CHAR_n  L500_CHAR_n_0
timestamp 1534323117
transform 1 0 224 0 1 136
box 0 0 12 18
use L500_CHAR_p  L500_CHAR_p_1
timestamp 1534323210
transform 1 0 240 0 1 136
box 0 0 12 18
use L500_CHAR_2  L500_CHAR_2_0
timestamp 1534324708
transform 1 0 256 0 1 136
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_CHAR_e  L500_CHAR_e_0
timestamp 1534321786
transform 1 0 114 0 1 50
box 0 0 12 18
use L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 173 0 1 50
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
