magic
tech scmos
timestamp 1542900940
use L500_CHAR_l  L500_CHAR_l_0 ../../Library/magic
timestamp 1534225390
transform 1 0 68 0 1 321
box 0 0 12 18
use L500_CHAR_i  L500_CHAR_i_0 ../../Library/magic
timestamp 1534226087
transform 1 0 84 0 1 321
box 0 0 8 18
use L500_CHAR_b  L500_CHAR_b_0 ../../Library/magic
timestamp 1534321628
transform 1 0 96 0 1 321
box 0 0 12 18
use L500_CHAR_r  L500_CHAR_r_0 ../../Library/magic
timestamp 1534323573
transform 1 0 112 0 1 321
box 0 0 12 18
use L500_CHAR_e  L500_CHAR_e_0 ../../Library/magic
timestamp 1534321786
transform 1 0 128 0 1 321
box 0 0 12 18
use L500_CHAR_s  L500_CHAR_s_0 ../../Library/magic
timestamp 1534323853
transform 1 0 148 0 1 321
box 0 0 12 18
use L500_CHAR_i  L500_CHAR_i_1
timestamp 1534226087
transform 1 0 164 0 1 321
box 0 0 8 18
use L500_CHAR_l  L500_CHAR_l_1
timestamp 1534225390
transform 1 0 176 0 1 321
box 0 0 12 18
use L500_CHAR_i  L500_CHAR_i_2
timestamp 1534226087
transform 1 0 192 0 1 321
box 0 0 8 18
use L500_CHAR_c  L500_CHAR_c_0 ../../Library/magic
timestamp 1534321654
transform 1 0 204 0 1 321
box 0 0 12 18
use L500_CHAR_o  L500_CHAR_o_0 ../../Library/magic
timestamp 1534323159
transform 1 0 220 0 1 321
box 0 0 12 18
use L500_CHAR_n  L500_CHAR_n_0 ../../Library/magic
timestamp 1534323117
transform 1 0 236 0 1 321
box 0 0 12 18
use T7_INV  T7_INV_0 ../../Library/magic
timestamp 1533657739
transform 1 0 32 0 1 163
box 0 0 16 56
use T11_NOR3  T11_NOR3_0 ../../Library/magic
timestamp 1533654861
transform 1 0 16 0 1 55
box 0 0 32 88
use L500_SIGNATURE_kallisti_big  L500_SIGNATURE_kallisti_big_0 ../../Library/magic
timestamp 1533657739
transform 1 0 45 0 1 67
box 9 8 231 235
use L500_SIGNATURE_pearlriver  L500_SIGNATURE_pearlriver_0 ../../Library/magic
timestamp 1542900699
transform 1 0 65 0 1 50
box 0 0 202 18
use T7_NAND2  T7_NAND2_0 ../../Library/magic
timestamp 1533654698
transform 0 1 24 -1 0 38
box 0 0 24 56
use T11_NOR2  T11_NOR2_0 ../../Library/magic
timestamp 1533654819
transform 0 1 86 -1 0 37
box 0 0 24 88
use T10_NAND2  T10_NAND2_0 ../../Library/magic
timestamp 1533654735
transform 0 1 179 -1 0 37
box 0 0 24 80
<< end >>
