magic
tech scmos
timestamp 1538814797
use Layout/magic/PearlRiver_quarter  PearlRiver_quarter_2
timestamp 1538814797
transform -1 0 7000 0 -1 8000
box 0 0 5900 3290
use Layout/magic/PearlRiver_quarter  PearlRiver_quarter_3
timestamp 1538814797
transform 0 1 2 -1 0 7000
box 0 0 5900 3290
use Layout/magic/PearlRiver_quarter  PearlRiver_quarter_1
timestamp 1538814797
transform 0 -1 8000 1 0 1000
box 0 0 5900 3290
use Layout/magic/PearlRiver_quarter  PearlRiver_quarter_0
timestamp 1538814797
transform 1 0 1000 0 1 0
box 0 0 5900 3290
<< end >>
