magic
tech scmos
timestamp 1540696282
<< error_s >>
rect 3252 2790 3254 3190
rect 3252 1364 3254 1370
rect 3252 1362 3274 1364
rect 3226 1322 3268 1324
rect 3272 1322 3274 1362
rect 3226 1318 3228 1322
rect 3232 1284 3234 1318
rect 3232 1282 3274 1284
rect 3226 1242 3268 1244
rect 3272 1242 3274 1282
rect 3226 1238 3228 1242
rect 3232 1204 3234 1238
rect 3232 1202 3274 1204
rect 3246 1162 3268 1164
rect 3272 1162 3274 1202
rect 3246 1158 3248 1162
rect 3252 1150 3254 1158
rect 2968 534 2992 539
rect 2994 534 3005 539
rect 2973 435 2974 534
rect 2987 435 2992 534
rect 2973 434 2992 435
rect 2999 435 3000 534
rect 3005 435 3010 534
rect 2999 434 3010 435
use Layout/magic/nmos_table  nmos_table_0
timestamp 1540696282
transform 1 0 750 0 1 850
box 0 0 1700 1700
use Layout/magic/metal1_rsquare  metal1_rsquare_0
timestamp 1540696282
transform 0 1 2500 1 0 850
box 0 0 2440 400
use diode_table  diode_table_0
timestamp 1540696282
transform 1 0 50 0 1 850
box 0 0 3104 2800
use Layout/magic/metal3_rsquare  metal3_rsquare_0
timestamp 1540696282
transform 0 1 2900 1 0 850
box 0 0 2440 400
use sonos_table  sonos_table_0
timestamp 1540696282
transform 1 0 -700 0 1 0
box 0 0 650 650
use Layout/magic/pad_measure  pad_measure_0
timestamp 1540696282
transform 0 1 0 -1 0 504
box 0 0 504 250
use Layout/magic/rpoly_rsquare  rpoly_rsquare_0
timestamp 1540696282
transform 1 0 300 0 1 400
box 0 0 2478 400
use hvnfet_table  hvnfet_table_0
timestamp 1540683310
transform 1 0 2852 0 1 407
box -3 -1 297 299
use Layout/magic/ringoscillator_stripe  ringoscillator_stripe_0
timestamp 1540696282
transform 0 1 3360 1 0 450
box 0 0 2704 440
use Layout/magic/pmos_table  pmos_table_0
timestamp 1540696282
transform 1 0 3900 0 1 450
box 0 0 1700 1700
use Layout/magic/caps_table  caps_table_0
timestamp 1540696282
transform 1 0 3900 0 1 450
box 0 0 2050 2072
use Layout/magic/polysi_rsquare  polysi_rsquare_0
timestamp 1540696282
transform 1 0 300 0 1 0
box 0 0 2478 400
use npn_table  npn_table_0
timestamp 1540696282
transform 1 0 2828 0 1 10
box 0 0 650 300
use Layout/magic/metal2_rsquare  metal2_rsquare_0
timestamp 1540696282
transform 1 0 3528 0 1 0
box 0 0 2440 400
<< end >>
