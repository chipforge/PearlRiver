magic
tech scmos
timestamp 1540699590
<< nwell >>
rect 110 180 190 190
rect 110 128 120 180
rect 131 156 169 169
rect 131 144 144 156
rect 156 144 169 156
rect 131 128 169 144
rect 180 128 190 180
rect 110 118 190 128
<< metal1 >>
rect 100 208 200 218
rect 145 178 155 208
rect 122 170 178 178
rect 122 130 130 170
rect 134 164 166 166
rect 134 160 136 164
rect 140 160 144 164
rect 148 160 152 164
rect 156 160 160 164
rect 164 160 166 164
rect 134 158 166 160
rect 134 156 142 158
rect 134 152 136 156
rect 140 152 142 156
rect 158 156 166 158
rect 134 148 142 152
rect 134 144 136 148
rect 140 144 142 148
rect 134 142 142 144
rect 146 85 154 154
rect 100 75 154 85
rect 158 152 160 156
rect 164 152 166 156
rect 158 148 166 152
rect 158 144 160 148
rect 164 144 166 148
rect 158 90 166 144
rect 170 130 178 170
rect 158 80 200 90
<< nwpbase >>
rect 120 169 180 180
rect 120 128 131 169
rect 144 144 156 156
rect 169 128 180 169
<< pbasepdiffcontact >>
rect 124 172 128 176
rect 132 172 136 176
rect 140 172 144 176
rect 148 172 152 176
rect 156 172 160 176
rect 164 172 168 176
rect 172 172 176 176
rect 124 164 128 168
rect 172 164 176 168
rect 124 156 128 160
rect 172 156 176 160
rect 124 148 128 152
rect 148 148 152 152
rect 172 148 176 152
rect 124 140 128 144
rect 172 140 176 144
rect 124 132 128 136
rect 172 132 176 136
<< nsubstratencontact >>
rect 136 160 140 164
rect 144 160 148 164
rect 152 160 156 164
rect 160 160 164 164
rect 136 152 140 156
rect 160 152 164 156
rect 136 144 140 148
rect 160 144 164 148
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_CHAR_c  L500_CHAR_c_0
timestamp 1534321654
transform 1 0 146 0 1 230
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_CHAR_p  L500_CHAR_p_0
timestamp 1534323117
transform 1 0 208 0 1 136
box 0 0 12 18
use L500_CHAR_n  L500_CHAR_n_0
timestamp 1534323210
transform 1 0 224 0 1 136
box 0 0 12 18
use L500_CHAR_p  L500_CHAR_p_1
timestamp 1534323117
transform 1 0 240 0 1 136
box 0 0 12 18
use L500_CHAR_1  L500_CHAR_1_0
timestamp 1534326485
transform 1 0 256 0 1 136
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_CHAR_e  L500_CHAR_e_0
timestamp 1534321786
transform 1 0 114 0 1 50
box 0 0 12 18
use L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 173 0 1 50
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
