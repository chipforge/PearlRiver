magic
tech scmos
timestamp 1540533428
<< polysilicon >>
rect 147 165 152 171
rect 147 131 152 137
<< metal1 >>
rect 90 181 100 200
rect 200 181 210 200
rect 90 171 145 181
rect 155 171 210 181
rect 90 121 145 131
rect 155 121 210 131
rect 90 100 100 121
rect 200 100 210 121
<< rndiffusion >>
rect 147 153 152 159
<< rpdiffusion >>
rect 147 143 152 149
<< rpoly >>
rect 147 149 152 153
<< polycontact >>
rect 145 171 155 181
rect 145 121 155 131
<< polyndiff >>
rect 147 159 152 165
<< polypdiff >>
rect 147 137 152 143
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
