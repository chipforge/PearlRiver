magic
tech scmos
timestamp 1534324363
<< metal1 >>
rect 0 14 4 18
rect 8 14 12 18
rect 0 12 12 14
rect 1 11 11 12
rect 3 10 9 11
rect 4 7 8 10
rect 3 6 9 7
rect 1 4 11 6
rect 0 3 12 4
rect 0 0 4 3
rect 8 0 12 3
<< end >>
