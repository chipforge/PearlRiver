magic
tech scmos
timestamp 1540530107
<< polysilicon >>
rect 140 165 160 177
rect 140 123 160 136
<< metal1 >>
rect 100 217 200 237
rect 140 197 160 217
rect 140 83 160 103
rect 100 63 200 83
<< rndiffusion >>
rect 140 152 160 165
<< rpdiffusion >>
rect 140 136 160 149
<< rpoly >>
rect 140 149 160 152
<< polycontact >>
rect 140 177 160 197
rect 140 103 160 123
use L500_TPAD_blank  L500_TPAD_blank_2 ./Library/magic
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
