magic
tech scmos
timestamp 1534325425
<< metal1 >>
rect 4 17 12 18
rect 2 16 12 17
rect 1 14 12 16
rect 0 13 6 14
rect 0 12 5 13
rect 0 4 4 12
rect 9 4 12 14
rect 0 0 12 4
<< end >>
