magic
tech scmos
timestamp 1534588197
<< metal1 >>
rect 2 17 10 18
rect 1 16 11 17
rect 0 14 12 16
rect 0 13 4 14
rect 8 13 12 14
rect 0 5 3 13
rect 9 7 12 13
rect 0 4 4 5
rect 7 4 12 7
rect 0 2 11 4
rect 1 1 11 2
rect 2 0 8 1
<< end >>
