magic
tech scmos
timestamp 1534323159
<< metal1 >>
rect 2 17 10 18
rect 1 16 11 17
rect 0 14 12 16
rect 0 4 4 14
rect 8 4 12 14
rect 0 2 12 4
rect 1 1 11 2
rect 2 0 10 1
<< end >>
