magic
tech scmos
timestamp 1534782471
<< nwell >>
rect 176 161 192 198
<< polysilicon >>
rect 175 179 179 181
rect 182 179 184 181
<< pdiffusion >>
rect 179 181 182 186
rect 179 173 182 179
<< metal1 >>
rect 90 224 100 248
rect 260 224 270 248
rect 90 214 146 224
rect 136 182 146 214
rect 178 214 270 224
rect 178 196 182 214
rect 136 178 165 182
rect 178 146 182 163
rect 90 136 182 146
rect 186 146 190 163
rect 186 136 270 146
rect 90 112 100 136
rect 260 112 270 136
<< ptransistor >>
rect 179 179 182 181
<< polycontact >>
rect 165 178 175 182
<< pdcontact >>
rect 178 186 182 196
rect 178 163 182 173
<< nsubstratencontact >>
rect 186 163 190 196
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_2 Library/magic
timestamp 1531942424
transform 1 0 0 0 1 240
box 0 0 120 120
use Library/magic/L500_CHAR_g  L500_CHAR_g_0 Library/magic
timestamp 1534322005
transform 1 0 120 0 1 230
box 0 0 12 18
use Library/magic/L500_CHAR_d  L500_CHAR_d_0 Library/magic
timestamp 1534321738
transform 1 0 228 0 1 230
box 0 0 12 18
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_3
timestamp 1531942424
transform 1 0 240 0 1 240
box 0 0 120 120
use Library/magic/L500_CHAR_3  L500_CHAR_3_0 Library/magic
timestamp 1534324785
transform 1 0 194 0 1 171
box 0 0 12 18
use Library/magic/L500_CHAR_slash  L500_CHAR_slash_0 Library/magic
timestamp 1534532558
transform 1 0 210 0 1 171
box 0 0 8 18
use Library/magic/L500_CHAR_2  L500_CHAR_2_1 Library/magic
timestamp 1534324708
transform 1 0 222 0 1 171
box 0 0 12 18
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_0
timestamp 1531942424
transform 1 0 0 0 1 0
box 0 0 120 120
use Library/magic/L500_CHAR_s  L500_CHAR_s_0 Library/magic
timestamp 1534323853
transform 1 0 120 0 1 112
box 0 0 12 18
use Library/magic/L500_CHAR_b  L500_CHAR_b_0 Library/magic
timestamp 1534321628
transform 1 0 228 0 1 112
box 0 0 12 18
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_1
timestamp 1531942424
transform 1 0 240 0 1 0
box 0 0 120 120
<< labels >>
rlabel space 20 260 100 340 1 gate
rlabel space 20 20 100 100 1 source
rlabel space 260 20 340 100 1 bulk
rlabel space 260 260 340 340 1 drain
<< end >>
