magic
tech scmos
timestamp 1541945102
<< nwell >>
rect 76 175 224 199
rect 76 125 100 175
rect 200 125 224 175
rect 76 101 224 125
<< metal1 >>
rect 83 192 217 200
rect 83 175 93 182
rect 207 175 217 182
rect 83 118 93 125
rect 107 129 193 132
rect 207 118 217 125
<< metal2 >>
rect 107 100 193 121
<< nwpbase >>
rect 100 125 200 175
<< pdcontact >>
rect 107 132 193 168
<< m2contact >>
rect 107 121 193 129
<< nsubstratencontact >>
rect 83 182 217 192
rect 83 125 93 175
rect 207 125 217 175
rect 83 108 217 118
use Library/magic/L500_CHAR_d  L500_CHAR_d_0 ~/IC/github/PearlRiver/Library/magic/Library/magic
timestamp 1534321738
transform 1 0 0 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_i  L500_CHAR_i_0 ~/IC/github/PearlRiver/Library/magic/Library/magic
timestamp 1534226087
transform 1 0 16 0 1 304
box 0 0 8 18
use Library/magic/L500_CHAR_o  L500_CHAR_o_1 ~/IC/github/PearlRiver/Library/magic/Library/magic
timestamp 1534323159
transform 1 0 28 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_d  L500_CHAR_d_1
timestamp 1534321738
transform 1 0 44 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_0 ~/IC/github/PearlRiver/Library/magic/Library/magic
timestamp 1534321786
transform 1 0 60 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_under  L500_CHAR_under_0 ~/IC/github/PearlRiver/Library/magic/Library/magic
timestamp 1534325915
transform 1 0 76 0 1 304
box 0 0 12 4
use Library/magic/L500_CHAR_p  L500_CHAR_p_0 ~/IC/github/PearlRiver/Library/magic/Library/magic
timestamp 1534323210
transform 1 0 92 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_b  L500_CHAR_b_0 ~/IC/github/PearlRiver/Library/magic/Library/magic
timestamp 1534321628
transform 1 0 108 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_0 Library/magic
timestamp 1534325357
transform 1 0 124 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_s  L500_CHAR_s_1 ~/IC/github/PearlRiver/Library/magic/Library/magic
timestamp 1534323853
transform 1 0 140 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_1
timestamp 1534321786
transform 1 0 156 0 1 304
box 0 0 12 18
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_0 Library/magic
timestamp 1537367970
transform 0 1 0 -1 0 300
box 0 0 100 300
use Library/magic/L500_CHAR_k  L500_CHAR_k_0 ~/IC/github/PearlRiver/Library/magic/Library/magic
timestamp 1534322894
transform 1 0 13 0 1 178
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_2
timestamp 1534325357
transform 1 0 225 0 1 141
box 0 0 12 18
use Library/magic/L500_CHAR_5  L500_CHAR_5_0 ~/IC/github/PearlRiver/Library/magic/Library/magic
timestamp 1534324893
transform 1 0 241 0 1 141
box 0 0 12 18
use Library/magic/L500_CHAR_tick  L500_CHAR_tick_0 ~/IC/github/PearlRiver/Library/magic/Library/magic
timestamp 1541212842
transform 1 0 257 0 1 141
box 0 12 4 18
use Library/magic/L500_CHAR_k  Library/magic/L500_CHAR_k_0
timestamp 1534322894
transform 1 0 265 0 1 141
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_1
timestamp 1534325357
transform 1 0 13 0 1 104
box 0 0 12 18
use Library/magic/L500_METAL2_W100_1rsquare  L500_METAL1_W100_2rsquare_0 Library/magic
timestamp 1537367970
transform 0 1 0 -1 0 100
box 0 0 100 300
<< end >>
