magic
tech scmos
timestamp 1531572553
<< nwell >>
rect 0 60 24 88
<< polysilicon >>
rect 7 78 9 80
rect 15 78 17 80
rect 7 60 9 62
rect 3 59 9 60
rect 6 58 9 59
rect 15 52 17 62
rect 15 51 21 52
rect 15 50 18 51
rect 6 17 9 18
rect 3 16 9 17
rect 7 14 9 16
rect 15 17 18 18
rect 15 16 21 17
rect 15 14 17 16
rect 7 8 9 10
rect 15 8 17 10
<< ndiffusion >>
rect 6 10 7 14
rect 9 10 10 14
rect 14 10 15 14
rect 17 10 18 14
<< pdiffusion >>
rect 6 62 7 78
rect 9 62 15 78
rect 17 62 18 78
<< metal1 >>
rect 2 78 6 82
rect 18 58 22 62
rect 2 30 6 55
rect 2 21 6 26
rect 10 54 22 58
rect 10 46 14 54
rect 10 14 14 42
rect 18 38 22 47
rect 18 21 22 34
rect 2 6 6 10
rect 18 6 22 10
<< ntransistor >>
rect 7 10 9 14
rect 15 10 17 14
<< ptransistor >>
rect 7 62 9 78
rect 15 62 17 78
<< polycontact >>
rect 2 55 6 59
rect 18 47 22 51
rect 2 17 6 21
rect 18 17 22 21
<< ndcontact >>
rect 2 10 6 14
rect 10 10 14 14
rect 18 10 22 14
<< pdcontact >>
rect 2 62 6 78
rect 18 62 22 78
<< m2contact >>
rect 2 26 6 30
rect 10 42 14 46
rect 18 34 22 38
<< psubstratepcontact >>
rect 0 2 24 6
<< nsubstratencontact >>
rect 0 82 24 86
<< labels >>
rlabel nsubstratencontact 2 82 24 86 5 vdd!
rlabel psubstratepcontact 2 2 24 6 1 gnd!
rlabel m2contact 2 26 6 30 3 B
rlabel m2contact 18 34 22 38 1 A
rlabel m2contact 10 42 14 46 1 Z
<< end >>
