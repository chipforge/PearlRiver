magic
tech scmos
timestamp 1542624506
<< nwell >>
rect 133 169 184 179
rect 133 130 143 169
rect 174 130 184 169
rect 133 120 184 130
<< pbasepolysilicon >>
rect 143 148 148 151
rect 156 148 159 151
<< metal1 >>
rect 100 200 143 210
rect 133 153 143 200
rect 200 164 210 200
rect 157 154 210 164
rect 90 135 148 145
rect 90 100 100 135
rect 162 100 172 135
rect 162 90 200 100
<< ntransistor >>
rect 148 148 156 151
<< nwpbase >>
rect 143 130 174 169
<< pbasendiffusion >>
rect 148 151 156 154
rect 148 145 156 148
<< pbasendiffcontact >>
rect 148 154 157 164
rect 148 135 157 145
<< pbasepdiffcontact >>
rect 162 135 172 151
<< polycontact >>
rect 133 148 143 153
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_CHAR_g  L500_CHAR_g_0
timestamp 1534322005
transform 1 0 101 0 1 178
box 0 0 12 18
use L500_CHAR_d  L500_CHAR_d_0
timestamp 1534321738
transform 1 0 184 0 1 187
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_CHAR_n  L500_CHAR_n_0
timestamp 1534323117
transform 1 0 215 0 1 140
box 0 0 12 18
use L500_CHAR_w  L500_CHAR_w_0
timestamp 1534324213
transform 1 0 235 0 1 152
box 0 0 16 18
use L500_CHAR_8  L500_CHAR_8_0
timestamp 1534324785
transform 1 0 255 0 1 152
box 0 0 12 18
use L500_CHAR_slash  L500_CHAR_slash_0
timestamp 1534532558
transform 1 0 271 0 1 152
box 0 0 8 18
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_CHAR_s  L500_CHAR_s_0
timestamp 1534323853
transform 1 0 104 0 1 95
box 0 0 12 18
use L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 190 0 1 104
box 0 0 12 18
use L500_CHAR_i  L500_CHAR_i_0
timestamp 1534226087
transform 1 0 215 0 1 118
box 0 0 8 18
use L500_CHAR_l  L500_CHAR_l_0
timestamp 1534225390
transform 1 0 239 0 1 130
box 0 0 12 18
use L500_CHAR_3  L500_CHAR_3_1
timestamp 1534324708
transform 1 0 255 0 1 130
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
