magic
tech scmos
timestamp 1539786992
<< polysilicon >>
rect 140 165 160 177
rect 140 123 160 135
<< metal1 >>
rect 80 197 100 200
rect 200 197 220 200
rect 80 177 140 197
rect 160 177 220 197
rect 80 103 140 123
rect 160 103 220 123
rect 80 100 100 103
rect 200 100 220 103
<< rndiffusion >>
rect 140 153 160 165
<< rpdiffusion >>
rect 140 135 160 147
<< rpoly >>
rect 140 147 160 153
<< polycontact >>
rect 140 177 160 197
rect 140 103 160 123
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
