magic
tech scmos
timestamp 1534325833
<< metal1 >>
rect 4 12 8 16
rect 0 8 12 12
rect 4 4 8 8
<< end >>
