magic
tech scmos
timestamp 1537375458
use Library/magic/L500_METAL1_W10_100rsquare  L500_METAL1_W10_100rsquare_0
timestamp 1537368500
transform 1 0 0 0 1 200
box 0 0 1200 100
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_1 Library/magic
timestamp 1537367970
transform 0 1 1100 -1 0 300
box 0 0 100 300
use Library/magic/L500_METAL1_W6_100rsquare  L500_METAL1_W6_100rsquare_0 Library/magic
timestamp 1537368500
transform 1 0 1300 0 1 200
box 0 0 800 100
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_2
timestamp 1537367970
transform 0 1 2000 -1 0 300
box 0 0 100 300
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_0
timestamp 1537367970
transform 1 0 0 0 1 0
box 0 0 100 300
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_4
timestamp 1537367970
transform 0 1 200 -1 0 180
box 0 0 100 300
use Library/magic/L500_METAL1_W8m_100rsquare  L500_METAL1_W8m_100rsquare_0
timestamp 1537373212
transform 1 0 400 0 1 80
box 0 0 640 100
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_5
timestamp 1537367970
transform 0 1 940 -1 0 180
box 0 0 100 300
use Library/magic/L500_METAL1_W4m_100rsquare  L500_METAL1_W4m_100rsquare_0
timestamp 1537372519
transform 1 0 1140 0 1 80
box 0 0 420 100
use Library/magic/L500_METAL1_W4_100rsquare  L500_METAL1_W4_100rsquare_0 Library/magic
timestamp 1537368500
transform 1 0 1460 0 1 80
box 0 0 600 100
use Library/magic/L500_METAL1_W20_100rsquare  L500_METAL1_W20_100rsquare_0 Library/magic
timestamp 1537368500
transform 1 0 0 0 1 0
box 0 0 2200 100
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_3
timestamp 1537367970
transform 0 1 2100 -1 0 100
box 0 0 100 300
use Library/magic/L500_METAL2_W100_1rsquare  L500_METAL2_W100_1rsquare_0 Library/magic
timestamp 1537367970
transform 1 0 1959 0 1 -120
box 0 0 100 300
<< end >>
