magic
tech scmos
timestamp 1534794778
use Layout/magic/L500_NMOS_table  L500_NMOS_table_0
timestamp 1534793986
transform 1 0 720 0 1 960
box 0 0 2280 2280
use Layout/magic/L500_RINGOSCILLATOR_stripe  L500_RINGOSCILLATOR_stripe_0
timestamp 1534793986
transform 0 1 3204 -1 0 3944
box 0 -114 2984 582
use Layout/magic/L500_PMOS_table  L500_PMOS_table_0 Layout/magic
timestamp 1534782471
transform 1 0 3880 0 1 960
box 0 0 2280 2280
use Layout/magic/L500_MOSFET_aligning  L500_MOSFET_aligning_0
timestamp 1533916061
transform 1 0 0 0 1 0
box 0 0 600 600
use Layout/magic/L500_METAL1_rsquare  L500_METAL1_rsquare_0
timestamp 1534793986
transform 1 0 720 0 1 480
box 0 0 2648 360
use Layout/magic/L500_METAL3_rsquare  L500_METAL3_rsquare_0
timestamp 1534793986
transform 1 0 3488 0 1 480
box 0 0 2532 360
use Layout/magic/L500_METAL2_rsquare  L500_METAL2_rsquare_0
timestamp 1534793986
transform 1 0 720 0 1 0
box 0 0 2648 360
use Layout/magic/L500_POLYSI_rsquare  L500_POLYSI_rsquare_0
timestamp 1534793986
transform 1 0 3488 0 1 0
box 0 0 2648 360
<< end >>
