magic
tech scmos
timestamp 1542621920
use L500_ZENER_W40_L1  L500_ZENER_W40_L1_0 ../../Library/magic
timestamp 1542620489
transform 1 0 2100 0 1 2100
box 0 0 304 300
use L500_ZENER_W40_L2  L500_ZENER_W40_L2_0 ../../Library/magic
timestamp 1542620489
transform 1 0 2450 0 1 2100
box 0 0 304 300
use L500_ZENER_W40_L3  L500_ZENER_W40_L3_0 ../../Library/magic
timestamp 1542620489
transform 1 0 2800 0 1 2100
box 0 0 304 300
use L500_ZENER_W40_L4  L500_ZENER_W40_L4_0 ../../Library/magic
timestamp 1542620489
transform 1 0 3150 0 1 2100
box 0 0 304 300
use L500_ZENER_W40_L5  L500_ZENER_W40_L5_0 ../../Library/magic
timestamp 1542620489
transform 1 0 3500 0 1 2100
box 0 0 304 300
use L500_ZENER_W20_L1  L500_ZENER_W20_L1_0 ../../Library/magic
timestamp 1540544127
transform 1 0 1750 0 1 1750
box 0 0 304 300
use L500_ZENER_W20_L2  L500_ZENER_W20_L2_0 ../../Library/magic
timestamp 1540543980
transform 1 0 2100 0 1 1750
box 0 0 304 300
use L500_ZENER_W20_L3  L500_ZENER_W20_L3_0 ../../Library/magic
timestamp 1540543901
transform 1 0 2450 0 1 1750
box 0 0 304 300
use L500_ZENER_W20_L4  L500_ZENER_W20_L4_0 ../../Library/magic
timestamp 1542620489
transform 1 0 2800 0 1 1750
box 0 0 304 300
use L500_ZENER_W20_L5  L500_ZENER_W20_L5_0 ../../Library/magic
timestamp 1540543671
transform 1 0 3150 0 1 1750
box 0 0 304 300
use L500_ZENER_W10_L5  L500_ZENER_W10_L5_0 ../../Library/magic
timestamp 1540543606
transform 1 0 1400 0 1 1400
box 0 0 304 300
use L500_ZENER_W5_L5  L500_ZENER_W5_L5_0 ../../Library/magic
timestamp 1540544708
transform 1 0 1750 0 1 1400
box 0 0 300 300
use L500_ZENER_W10_L4  L500_ZENER_W10_L4_0 ../../Library/magic
timestamp 1542620489
transform 1 0 1050 0 1 1050
box 0 0 304 300
use L500_ZENER_W5_L4  L500_ZENER_W5_L4_0 ../../Library/magic
timestamp 1542620489
transform 1 0 1400 0 1 1050
box 0 0 300 300
use L500_DIODE_PBASE_A2k_params  L500_DIODE_PBASE_A2k_params_0 ../../Library/magic
timestamp 1541945167
transform 1 0 3152 0 1 1299
box 0 0 300 322
use L500_DIODE_PBASE_A10k_params  L500_DIODE_PBASE_A10k_params_0 ../../Library/magic
timestamp 1541995960
transform 1 0 3498 0 1 1299
box 0 0 301 322
use L500_ZENER_W10_L3  L500_ZENER_W10_L3_0 ../../Library/magic
timestamp 1540543464
transform 1 0 700 0 1 700
box 0 0 304 300
use L500_ZENER_W5_L3  L500_ZENER_W5_L3_0 ../../Library/magic
timestamp 1540544786
transform 1 0 1050 0 1 700
box 0 0 300 300
use L500_DIODE_SUBSTRATE_A1k_params  L500_DIODE_SUBSTRATE_A1k_params_0 ../../Library/magic
timestamp 1541215827
transform 1 0 3152 0 1 949
box 0 0 300 322
use L500_DIODE_SUBSTRATE_A10k_params  L500_DIODE_SUBSTRATE_A10k_params_0 ../../Library/magic
timestamp 1541224905
transform 1 0 3498 0 1 949
box 0 0 301 322
use L500_ZENER_W10_L2  L500_ZENER_W10_L2_0 ../../Library/magic
timestamp 1540542704
transform 1 0 350 0 1 350
box 0 0 304 300
use L500_ZENER_W5_L2  L500_ZENER_W5_L2_0 ../../Library/magic
timestamp 1540544905
transform 1 0 700 0 1 350
box 0 0 300 300
use L500_ZENER_W10_L1  L500_ZENER_W10_L1_0 ../../Library/magic
timestamp 1540539143
transform 1 0 0 0 1 0
box 0 0 304 300
use L500_ZENER_W5_L1  L500_ZENER_W5_L1_0 ../../Library/magic
timestamp 1540544919
transform 1 0 350 0 1 0
box 0 0 300 300
<< end >>
