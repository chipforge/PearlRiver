magic
tech scmos
timestamp 1534325915
<< metal1 >>
rect 0 0 12 4
<< end >>
