magic
tech scmos
timestamp 1540531615
<< polysilicon >>
rect 147 159 152 165
rect 147 134 152 140
<< metal1 >>
rect 90 175 100 200
rect 200 175 210 200
rect 90 165 145 175
rect 155 165 210 175
rect 90 124 145 134
rect 155 124 210 134
rect 90 100 100 124
rect 200 100 210 124
<< rndiffusion >>
rect 147 150 152 153
<< rpdiffusion >>
rect 147 146 152 149
<< rpoly >>
rect 147 149 152 150
<< polycontact >>
rect 145 165 155 175
rect 145 124 155 134
<< polyndiff >>
rect 147 153 152 159
<< polypdiff >>
rect 147 140 152 146
use L500_TPAD_blank  L500_TPAD_blank_2 ./Library/magic
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
