magic
tech scmos
timestamp 1540616762
use Library/magic/L500_ZENER_W5_L5  L500_ZENER_W5_L5_0
timestamp 1540544708
transform 1 0 1750 0 1 1400
box 0 0 300 300
use Library/magic/L500_ZENER_W5_L4  L500_ZENER_W5_L4_0
timestamp 1540544728
transform 1 0 1400 0 1 1050
box 0 0 300 300
use Library/magic/L500_ZENER_W5_L3  L500_ZENER_W5_L3_0
timestamp 1540544786
transform 1 0 1050 0 1 700
box 0 0 300 300
use Library/magic/L500_ZENER_W5_L2  L500_ZENER_W5_L2_0
timestamp 1540544905
transform 1 0 700 0 1 350
box 0 0 300 300
use Library/magic/L500_ZENER_W5_L1  L500_ZENER_W5_L1_0
timestamp 1540544919
transform 1 0 350 0 1 0
box 0 0 300 300
use Library/magic/L500_ZENER_W10_L5  L500_ZENER_W10_L5_0
timestamp 1540544708
transform 1 0 1400 0 1 1400
box 0 0 300 300
use Library/magic/L500_ZENER_W10_L4  L500_ZENER_W10_L4_0
timestamp 1540544728
transform 1 0 1050 0 1 1050
box 0 0 300 300
use Library/magic/L500_ZENER_W10_L3  L500_ZENER_W10_L3_0
timestamp 1540544786
transform 1 0 700 0 1 700
box 0 0 300 300
use Library/magic/L500_ZENER_W10_L2  L500_ZENER_W10_L2_0
timestamp 1540544905
transform 1 0 350 0 1 350 
box 0 0 300 300
use Library/magic/L500_ZENER_W10_L1  L500_ZENER_W10_L1_0
timestamp 1540544919
transform 1 0 0 0 1 0 
box 0 0 300 300
use Library/magic/L500_ZENER_W20_L1  L500_ZENER_W20_L1_0
timestamp 1540544708
transform 1 0 1750 0 1 1750
box 0 0 300 300
use Library/magic/L500_ZENER_W20_L2  L500_ZENER_W20_L2_0
timestamp 1540544708
transform 1 0 2100 0 1 1750
box 0 0 300 300
use Library/magic/L500_ZENER_W20_L3  L500_ZENER_W20_L3_0
timestamp 1540544708
transform 1 0 2450 0 1 1750
box 0 0 300 300
use Library/magic/L500_ZENER_W20_L4  L500_ZENER_W20_L4_0
timestamp 1540544708
transform 1 0 2800 0 1 1750
box 0 0 300 300
use Library/magic/L500_ZENER_W20_L5  L500_ZENER_W20_L5_0
timestamp 1540544708
transform 1 0 3150 0 1 1750
box 0 0 300 300
use Library/magic/L500_ZENER_W40_L1  L500_ZENER_W40_L1_0
timestamp 1540544708
transform 1 0 2100 0 1 2100
box 0 0 300 300
use Library/magic/L500_ZENER_W40_L2  L500_ZENER_W40_L2_0
timestamp 1540544708
transform 1 0 2450 0 1 2100
box 0 0 300 300
use Library/magic/L500_ZENER_W40_L3  L500_ZENER_W40_L3_0
timestamp 1540544708
transform 1 0 2800 0 1 2100
box 0 0 300 300
use Library/magic/L500_ZENER_W40_L4  L500_ZENER_W40_L4_0
timestamp 1540544708
transform 1 0 3150 0 1 2100
box 0 0 300 300
use Library/magic/L500_ZENER_W40_L5  L500_ZENER_W40_L5_0
timestamp 1540544708
transform 1 0 3500 0 1 2100
box 0 0 300 300
<< end >>
