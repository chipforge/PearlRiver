magic
tech scmos
timestamp 1531683380
<< nwell >>
rect 0 58 32 88
<< polysilicon >>
rect 7 78 9 80
rect 12 78 14 80
rect 17 78 19 80
rect 7 58 9 60
rect 3 57 9 58
rect 6 56 9 57
rect 12 54 14 60
rect 17 58 19 60
rect 17 57 21 58
rect 17 56 18 57
rect 12 53 15 54
rect 14 50 15 53
rect 14 25 15 28
rect 22 25 23 28
rect 13 22 15 25
rect 21 22 23 25
rect 13 20 17 22
rect 21 20 25 22
rect 6 17 9 18
rect 3 16 9 17
rect 7 13 9 16
rect 15 13 17 20
rect 23 13 25 20
rect 7 8 9 10
rect 15 8 17 10
rect 23 8 25 10
<< ndiffusion >>
rect 6 10 7 13
rect 9 10 10 13
rect 14 10 15 13
rect 17 10 18 13
rect 22 10 23 13
rect 25 10 26 13
<< pdiffusion >>
rect 6 60 7 78
rect 9 60 12 78
rect 14 60 17 78
rect 19 60 20 78
<< metal1 >>
rect 30 82 32 86
rect 2 78 6 82
rect 25 60 30 64
rect 2 30 6 53
rect 2 21 6 26
rect 10 46 14 49
rect 10 29 14 42
rect 18 38 22 53
rect 18 29 22 34
rect 26 54 30 60
rect 26 22 30 50
rect 10 18 26 22
rect 10 14 14 18
rect 26 14 30 18
rect 2 6 6 10
rect 18 6 22 10
rect 30 2 32 6
<< metal2 >>
rect 2 82 30 86
rect 2 2 30 6
<< ntransistor >>
rect 7 10 9 13
rect 15 10 17 13
rect 23 10 25 13
<< ptransistor >>
rect 7 60 9 78
rect 12 60 14 78
rect 17 60 19 78
<< polycontact >>
rect 2 53 6 57
rect 18 53 22 57
rect 10 49 14 53
rect 10 25 14 29
rect 18 25 22 29
rect 2 17 6 21
<< ndcontact >>
rect 2 10 6 14
rect 10 10 14 14
rect 18 10 22 14
rect 26 10 30 14
<< pdcontact >>
rect 2 60 6 78
rect 20 60 25 78
<< m2contact >>
rect 2 26 6 30
rect 10 42 14 46
rect 18 34 22 38
rect 26 50 30 54
rect 26 18 30 22
<< psubstratepcontact >>
rect 0 2 30 6
<< nsubstratencontact >>
rect 0 82 30 86
<< labels >>
rlabel nsubstratencontact 2 82 30 86 5 vdd!
rlabel psubstratepcontact 2 2 30 6 1 gnd!
rlabel m2contact 18 34 22 38 1 A
rlabel m2contact 26 50 30 54 1 Z
rlabel m2contact 10 42 14 46 1 B
rlabel m2contact 2 26 6 30 3 C
rlabel m2contact 26 18 30 22 7 Z
<< end >>
