magic
tech scmos
timestamp 1534326416
<< error_s >>
rect 192 18 197 19
use Library/magic/L500_CHAR_p  L500_CHAR_p_0 Library/magic
timestamp 1534323210
transform 1 0 0 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_0 Library/magic
timestamp 1534321786
transform 1 0 16 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_0 Library/magic
timestamp 1534325357
transform 1 0 32 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_r  L500_CHAR_r_0 Library/magic
timestamp 1534323573
transform 1 0 48 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_l  L500_CHAR_l_0 Library/magic
timestamp 1534225390
transform 1 0 64 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_r  L500_CHAR_r_1
timestamp 1534323573
transform 1 0 80 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_i  L500_CHAR_i_0 Library/magic
timestamp 1534226087
transform 1 0 96 0 1 0
box 0 0 8 18
use Library/magic/L500_CHAR_v  L500_CHAR_v_0 Library/magic
timestamp 1534324131
transform 1 0 108 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_1
timestamp 1534321786
transform 1 0 124 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_r  L500_CHAR_r_2
timestamp 1534323573
transform 1 0 140 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_v  L500_CHAR_v_1
timestamp 1534324131
transform 1 0 168 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_dot  L500_CHAR_dot_0 Library/magic
timestamp 1534325697
transform 1 0 182 0 1 0
box 0 0 4 4
use Library/magic/L500_CHAR_1  L500_CHAR_1_0 Library/magic
timestamp 1534319458
transform 1 0 190 0 1 0
box 0 0 12 18
<< end >>
