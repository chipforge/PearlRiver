magic
tech scmos
timestamp 1534324893
<< metal1 >>
rect 0 15 12 18
rect 0 11 4 15
rect 0 10 10 11
rect 0 9 11 10
rect 0 8 12 9
rect 7 7 12 8
rect 8 4 12 7
rect 0 2 12 4
rect 0 1 11 2
rect 0 0 10 1
<< end >>
