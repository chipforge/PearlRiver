magic
tech scmos
timestamp 1534782471
<< metal1 >>
rect -352 152 0 156
rect 824 152 1176 156
rect -352 135 -328 152
rect -316 135 -304 152
rect -294 135 -284 152
rect -276 135 -268 152
rect -262 135 -256 152
rect -252 135 -248 152
rect 1072 130 1076 152
rect 1080 130 1086 152
rect 1092 130 1100 152
rect 1108 130 1118 152
rect 1128 130 1140 152
rect 1152 130 1176 152
rect -8 80 0 84
rect 824 80 832 84
rect -8 72 0 76
rect 824 72 832 76
rect -352 4 -348 32
rect -344 4 -338 32
rect -332 4 -324 32
rect -316 4 -306 32
rect -296 4 -284 32
rect -272 4 -248 32
rect 1072 4 1076 32
rect 1080 4 1086 32
rect 1092 4 1100 32
rect 1108 4 1118 32
rect 1128 4 1140 32
rect 1152 4 1176 32
rect -352 0 19 4
rect 824 0 1176 4
<< metal2 >>
rect 810 128 814 164
rect 18 116 22 124
rect 50 116 54 124
rect 82 116 86 124
rect 114 116 118 124
rect 146 116 150 124
rect 178 116 182 124
rect 210 116 214 124
rect 242 116 246 124
rect 274 116 278 124
rect 306 116 310 124
rect 338 116 342 124
rect 370 116 374 124
rect 402 116 406 124
rect 434 116 438 124
rect 466 116 470 124
rect 498 116 502 124
rect 530 116 534 124
rect 562 116 566 124
rect 594 116 598 124
rect 626 116 630 124
rect 658 116 662 124
rect 690 116 694 124
rect 722 116 726 124
rect 754 116 758 124
rect 786 116 790 124
rect 802 116 806 124
rect 10 112 30 116
rect 42 112 62 116
rect 74 112 94 116
rect 106 112 126 116
rect 138 112 158 116
rect 170 112 190 116
rect 202 112 222 116
rect 234 112 254 116
rect 266 112 286 116
rect 298 112 318 116
rect 330 112 350 116
rect 362 112 382 116
rect 394 112 414 116
rect 426 112 446 116
rect 458 112 478 116
rect 490 112 510 116
rect 522 112 542 116
rect 554 112 574 116
rect 586 112 606 116
rect 618 112 638 116
rect 650 112 670 116
rect 682 112 702 116
rect 714 112 734 116
rect 746 112 766 116
rect 778 112 818 116
rect 26 108 30 112
rect 58 108 62 112
rect 90 108 94 112
rect 122 108 126 112
rect 154 108 158 112
rect 186 108 190 112
rect 218 108 222 112
rect 250 108 254 112
rect 282 108 286 112
rect 314 108 318 112
rect 346 108 350 112
rect 378 108 382 112
rect 410 108 414 112
rect 442 108 446 112
rect 474 108 478 112
rect 506 108 510 112
rect 538 108 542 112
rect 570 108 574 112
rect 602 108 606 112
rect 634 108 638 112
rect 666 108 670 112
rect 698 108 702 112
rect 730 108 734 112
rect 762 108 766 112
rect 26 104 38 108
rect 58 104 70 108
rect 90 104 102 108
rect 122 104 134 108
rect 154 104 166 108
rect 186 104 198 108
rect 218 104 230 108
rect 250 104 262 108
rect 282 104 294 108
rect 314 104 326 108
rect 346 104 358 108
rect 378 104 390 108
rect 410 104 422 108
rect 442 104 454 108
rect 474 104 486 108
rect 506 104 518 108
rect 538 104 550 108
rect 570 104 582 108
rect 602 104 614 108
rect 634 104 646 108
rect 666 104 678 108
rect 698 104 710 108
rect 730 104 742 108
rect 762 104 774 108
rect 2 40 6 100
rect 34 96 38 104
rect 66 96 70 104
rect 98 96 102 104
rect 130 96 134 104
rect 162 96 166 104
rect 194 96 198 104
rect 226 96 230 104
rect 258 96 262 104
rect 290 96 294 104
rect 322 96 326 104
rect 354 96 358 104
rect 386 96 390 104
rect 418 96 422 104
rect 450 96 454 104
rect 482 96 486 104
rect 514 96 518 104
rect 546 96 550 104
rect 578 96 582 104
rect 610 96 614 104
rect 642 96 646 104
rect 674 96 678 104
rect 706 96 710 104
rect 738 96 742 104
rect 770 96 774 104
rect 794 100 798 112
rect 794 96 806 100
rect 802 60 806 96
rect 50 52 54 60
rect 82 52 86 60
rect 114 52 118 60
rect 146 52 150 60
rect 178 52 182 60
rect 210 52 214 60
rect 242 52 246 60
rect 274 52 278 60
rect 306 52 310 60
rect 338 52 342 60
rect 370 52 374 60
rect 402 52 406 60
rect 434 52 438 60
rect 466 52 470 60
rect 498 52 502 60
rect 530 52 534 60
rect 562 52 566 60
rect 594 52 598 60
rect 626 52 630 60
rect 658 52 662 60
rect 690 52 694 60
rect 722 52 726 60
rect 754 52 758 60
rect 786 52 790 60
rect 802 56 822 60
rect 10 48 30 52
rect 50 48 62 52
rect 82 48 94 52
rect 114 48 126 52
rect 146 48 158 52
rect 178 48 190 52
rect 210 48 222 52
rect 242 48 254 52
rect 274 48 286 52
rect 306 48 318 52
rect 338 48 350 52
rect 370 48 382 52
rect 402 48 414 52
rect 434 48 446 52
rect 466 48 478 52
rect 498 48 510 52
rect 530 48 542 52
rect 562 48 574 52
rect 594 48 606 52
rect 626 48 638 52
rect 658 48 670 52
rect 690 48 702 52
rect 722 48 734 52
rect 754 48 766 52
rect 786 48 798 52
rect 26 44 30 48
rect 58 44 62 48
rect 90 44 94 48
rect 122 44 126 48
rect 154 44 158 48
rect 186 44 190 48
rect 218 44 222 48
rect 250 44 254 48
rect 282 44 286 48
rect 314 44 318 48
rect 346 44 350 48
rect 378 44 382 48
rect 410 44 414 48
rect 442 44 446 48
rect 474 44 478 48
rect 506 44 510 48
rect 538 44 542 48
rect 570 44 574 48
rect 602 44 606 48
rect 634 44 638 48
rect 666 44 670 48
rect 698 44 702 48
rect 730 44 734 48
rect 762 44 766 48
rect 794 44 798 48
rect 26 40 46 44
rect 58 40 78 44
rect 90 40 110 44
rect 122 40 142 44
rect 154 40 174 44
rect 186 40 206 44
rect 218 40 238 44
rect 250 40 270 44
rect 282 40 302 44
rect 314 40 334 44
rect 346 40 366 44
rect 378 40 398 44
rect 410 40 430 44
rect 442 40 462 44
rect 474 40 494 44
rect 506 40 526 44
rect 538 40 558 44
rect 570 40 590 44
rect 602 40 622 44
rect 634 40 654 44
rect 666 40 686 44
rect 698 40 718 44
rect 730 40 750 44
rect 762 40 782 44
rect 794 40 814 44
rect 18 -8 22 36
rect 34 32 38 40
rect 66 32 70 40
rect 98 32 102 40
rect 130 32 134 40
rect 162 32 166 40
rect 194 32 198 40
rect 226 32 230 40
rect 258 32 262 40
rect 290 32 294 40
rect 322 32 326 40
rect 354 32 358 40
rect 386 32 390 40
rect 418 32 422 40
rect 450 32 454 40
rect 482 32 486 40
rect 514 32 518 40
rect 546 32 550 40
rect 578 32 582 40
rect 610 32 614 40
rect 642 32 646 40
rect 674 32 678 40
rect 706 32 710 40
rect 738 32 742 40
rect 770 32 774 40
rect 802 32 806 40
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_1 Library/magic
timestamp 1531942424
transform 1 0 -360 0 1 24
box 0 0 120 120
use Library/magic/L500_SIGNATURE_vdd  L500_SIGNATURE_vdd_0 Library/magic
timestamp 1534327146
transform 1 0 -172 0 1 100
box 0 0 52 18
use Library/magic/L500_SIGNATURE_gnd  L500_SIGNATURE_gnd_0 Library/magic
timestamp 1534327291
transform 1 0 -240 0 1 38
box 0 0 52 18
use Library/magic/T10_NAND3  T10_NAND3_49 Library/magic
timestamp 1533654785
transform -1 0 32 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_48
timestamp 1533654785
transform -1 0 64 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_47
timestamp 1533654785
transform -1 0 96 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_46
timestamp 1533654785
transform -1 0 128 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_45
timestamp 1533654785
transform -1 0 160 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_44
timestamp 1533654785
transform -1 0 192 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_43
timestamp 1533654785
transform -1 0 224 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_42
timestamp 1533654785
transform -1 0 256 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_41
timestamp 1533654785
transform -1 0 288 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_40
timestamp 1533654785
transform -1 0 320 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_39
timestamp 1533654785
transform -1 0 352 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_38
timestamp 1533654785
transform -1 0 384 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_37
timestamp 1533654785
transform -1 0 416 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_36
timestamp 1533654785
transform -1 0 448 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_35
timestamp 1533654785
transform -1 0 480 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_34
timestamp 1533654785
transform -1 0 512 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_33
timestamp 1533654785
transform -1 0 544 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_32
timestamp 1533654785
transform -1 0 576 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_31
timestamp 1533654785
transform -1 0 608 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_30
timestamp 1533654785
transform -1 0 640 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_29
timestamp 1533654785
transform -1 0 672 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_28
timestamp 1533654785
transform -1 0 704 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_27
timestamp 1533654785
transform -1 0 736 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_26
timestamp 1533654785
transform -1 0 768 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_25
timestamp 1533654785
transform -1 0 800 0 -1 158
box 0 0 32 80
use Library/magic/T10_NAND2  T10_NAND2_1 Library/magic
timestamp 1533654735
transform -1 0 824 0 -1 158
box 0 0 24 80
use Library/magic/L500_CHAR_r  L500_CHAR_r_0 Library/magic
timestamp 1534323573
transform 1 0 -240 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_o  L500_CHAR_o_0 Library/magic
timestamp 1534323159
transform 1 0 -224 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_5  L500_CHAR_5_0 Library/magic
timestamp 1534324893
transform 1 0 -208 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_1  L500_CHAR_1_0 Library/magic
timestamp 1534326485
transform 1 0 -192 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_under  L500_CHAR_under_0 Library/magic
timestamp 1534325915
transform 1 0 -176 0 1 8
box 0 0 12 4
use Library/magic/L500_CHAR_n  L500_CHAR_n_0 Library/magic
timestamp 1534323117
transform 1 0 -160 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_0 Library/magic
timestamp 1534325357
transform 1 0 -144 0 1 8
box 0 0 12 18
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_0
timestamp 1531942424
transform 1 0 -120 0 1 24
box 0 0 120 120
use Library/magic/L500_CHAR_n  L500_CHAR_n_1
timestamp 1534323117
transform 1 0 -128 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_d  L500_CHAR_d_0 Library/magic
timestamp 1534321738
transform 1 0 -112 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_3  L500_CHAR_3_0 Library/magic
timestamp 1534324785
transform 1 0 -96 0 1 8
box 0 0 12 18
use Library/magic/T10_NAND2  T10_NAND2_0
timestamp 1533654735
transform 1 0 0 0 1 -2
box 0 0 24 80
use Library/magic/T10_NAND3  T10_NAND3_0
timestamp 1533654785
transform 1 0 24 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_1
timestamp 1533654785
transform 1 0 56 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_2
timestamp 1533654785
transform 1 0 88 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_3
timestamp 1533654785
transform 1 0 120 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_4
timestamp 1533654785
transform 1 0 152 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_5
timestamp 1533654785
transform 1 0 184 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_6
timestamp 1533654785
transform 1 0 216 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_7
timestamp 1533654785
transform 1 0 248 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_8
timestamp 1533654785
transform 1 0 280 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_9
timestamp 1533654785
transform 1 0 312 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_10
timestamp 1533654785
transform 1 0 344 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_11
timestamp 1533654785
transform 1 0 376 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_12
timestamp 1533654785
transform 1 0 408 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_13
timestamp 1533654785
transform 1 0 440 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_14
timestamp 1533654785
transform 1 0 472 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_15
timestamp 1533654785
transform 1 0 504 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_16
timestamp 1533654785
transform 1 0 536 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_17
timestamp 1533654785
transform 1 0 568 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_18
timestamp 1533654785
transform 1 0 600 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_19
timestamp 1533654785
transform 1 0 632 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_20
timestamp 1533654785
transform 1 0 664 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_21
timestamp 1533654785
transform 1 0 696 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_22
timestamp 1533654785
transform 1 0 728 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_23
timestamp 1533654785
transform 1 0 760 0 1 -2
box 0 0 32 80
use Library/magic/T10_NAND3  T10_NAND3_24
timestamp 1533654785
transform 1 0 792 0 1 -2
box 0 0 32 80
use Library/magic/L500_SIGNATURE_vdd  L500_SIGNATURE_vdd_1
timestamp 1534327146
transform 1 0 944 0 1 100
box 0 0 52 18
use Library/magic/L500_SIGNATURE_gnd  L500_SIGNATURE_gnd_1
timestamp 1534327291
transform 1 0 1012 0 1 38
box 0 0 52 18
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_2
timestamp 1531942424
transform 1 0 824 0 1 24
box 0 0 120 120
use Library/magic/L500_CHAR_r  L500_CHAR_r_1
timestamp 1534323573
transform 1 0 908 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_o  L500_CHAR_o_1
timestamp 1534323159
transform 1 0 924 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_5  L500_CHAR_5_1
timestamp 1534324893
transform 1 0 940 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_1  L500_CHAR_1_1
timestamp 1534326485
transform 1 0 956 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_under  L500_CHAR_under_1
timestamp 1534325915
transform 1 0 972 0 1 8
box 0 0 12 4
use Library/magic/L500_CHAR_n  L500_CHAR_n_2
timestamp 1534323117
transform 1 0 988 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_1
timestamp 1534325357
transform 1 0 1004 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_n  L500_CHAR_n_3
timestamp 1534323117
transform 1 0 1020 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_d  L500_CHAR_d_1
timestamp 1534321738
transform 1 0 1036 0 1 8
box 0 0 12 18
use Library/magic/L500_CHAR_3  L500_CHAR_3_1
timestamp 1534324785
transform 1 0 1052 0 1 8
box 0 0 12 18
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_3
timestamp 1531942424
transform 1 0 1064 0 1 24
box 0 0 120 120
<< labels >>
rlabel space -100 44 -20 118 1 vdd!
rlabel space -340 44 -260 118 1 gnd!
rlabel space 844 44 924 118 1 vdd!
rlabel space 1084 44 1164 118 1 gnd!
rlabel metal2 18 -8 22 -4 1 en
rlabel metal2 810 160 814 164 5 out
<< end >>
