magic
tech scmos
timestamp 1534325697
<< metal1 >>
rect 0 0 4 4
<< end >>
