magic
tech scmos
timestamp 1534323899
<< metal1 >>
rect 0 4 4 18
rect 8 4 12 18
rect 0 1 12 4
rect 1 0 11 1
<< end >>
