magic
tech scmos
timestamp 1534323446
<< metal1 >>
rect 2 17 10 18
rect 1 16 11 17
rect 0 14 12 16
rect 0 5 4 14
rect 8 13 12 14
rect 9 7 12 13
rect 8 6 12 7
rect 8 5 13 6
rect 0 4 5 5
rect 8 4 14 5
rect 0 2 14 4
rect 1 1 13 2
rect 2 0 11 1
<< end >>
