magic
tech scmos
timestamp 1539444003
<< nwell >>
rect -6 -10 43 28
<< pbasepolysilicon >>
rect 16 18 20 22
rect 16 8 20 10
<< sonostransistor >>
rect 16 10 20 18
<< pbase >>
rect 0 18 16 22
rect 20 18 37 22
rect 0 10 4 18
rect 32 10 37 18
rect 0 8 16 10
rect 20 8 37 10
rect 0 4 37 8
rect 0 0 4 4
rect 32 0 37 4
rect 0 -4 37 0
<< polycontact >>
rect 16 22 20 26
<< pbasendiffusion >>
rect 12 10 16 18
rect 20 10 24 18
<< pbasendiffcontact >>
rect 4 10 12 18
rect 24 10 32 18
<< pbasepdiffcontact >>
rect 4 0 32 4
<< end >>
