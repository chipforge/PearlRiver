magic
tech scmos
timestamp 1538569292
<< metal2 >>
rect 1765 310 1773 314
rect 1769 292 1773 310
rect 2185 310 2204 314
rect 2185 295 2189 310
rect 300 274 308 278
rect 1120 274 1136 278
rect 300 178 308 182
rect 1120 178 1136 182
use Layout/magic/T10_RO51_NAND3  T10_RO51_NAND3_0
timestamp 1538561894
transform 1 0 310 0 -1 438
box -310 -2 1126 180
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_2 Library/magic
timestamp 1537343441
transform 1 0 1665 0 1 310
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 2204 0 1 310
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 200 0 1 178
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 1136 0 1 178
box 0 0 100 100
use Layout/magic/T11_RO51_NOR3  T11_RO51_NOR3_0
timestamp 1538561069
transform 1 0 310 0 1 2
box -310 -2 1126 196
use Layout/magic/T7_RO51_INV  T7_RO51_INV_0
timestamp 1538566008
transform 1 0 1775 0 1 169
box -310 -2 728 142
use Layout/magic/T7_CELL50_FILLCAP  T7_CELL50_FILLCAP_0
timestamp 1538559977
transform 1 0 2911 0 1 169
box -310 -2 904 140
<< end >>
