magic
tech scmos
timestamp 1534323853
<< metal1 >>
rect 2 17 12 18
rect 1 16 12 17
rect 0 15 12 16
rect 0 14 5 15
rect 9 14 12 15
rect 0 11 4 14
rect 0 10 6 11
rect 0 9 11 10
rect 1 8 12 9
rect 3 7 12 8
rect 8 4 12 7
rect 0 3 3 4
rect 6 3 12 4
rect 0 2 12 3
rect 0 1 11 2
rect 0 0 10 1
<< end >>
