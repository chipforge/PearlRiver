magic
tech scmos
timestamp 1540701346
<< nwell >>
rect 106 184 194 194
rect 106 124 116 184
rect 128 160 172 172
rect 128 140 140 160
rect 160 140 172 160
rect 128 124 172 140
rect 184 124 194 184
rect 106 114 194 124
<< metal1 >>
rect 100 208 200 218
rect 145 182 155 208
rect 118 174 182 182
rect 118 126 126 174
rect 130 168 170 170
rect 130 164 132 168
rect 136 164 140 168
rect 144 164 148 168
rect 152 164 156 168
rect 160 164 164 168
rect 168 164 170 168
rect 130 162 170 164
rect 130 160 138 162
rect 130 156 132 160
rect 136 156 138 160
rect 162 160 170 162
rect 130 152 138 156
rect 130 148 132 152
rect 136 148 138 152
rect 130 144 138 148
rect 130 140 132 144
rect 136 140 138 144
rect 130 136 138 140
rect 130 132 132 136
rect 136 132 138 136
rect 130 130 138 132
rect 142 142 158 158
rect 162 156 164 160
rect 168 156 170 160
rect 162 152 170 156
rect 162 148 164 152
rect 168 148 170 152
rect 162 144 170 148
rect 142 85 152 142
rect 100 75 152 85
rect 162 140 164 144
rect 168 140 170 144
rect 162 136 170 140
rect 162 132 164 136
rect 168 132 170 136
rect 162 90 170 132
rect 174 126 182 174
rect 162 80 200 90
<< nwpbase >>
rect 116 172 184 184
rect 116 124 128 172
rect 140 140 160 160
rect 172 124 184 172
<< pbasepdiffcontact >>
rect 120 176 124 180
rect 128 176 132 180
rect 136 176 140 180
rect 144 176 148 180
rect 152 176 156 180
rect 160 176 164 180
rect 168 176 172 180
rect 176 176 180 180
rect 120 168 124 172
rect 176 168 180 172
rect 120 160 124 164
rect 176 160 180 164
rect 120 152 124 156
rect 144 152 148 156
rect 152 152 156 156
rect 176 152 180 156
rect 120 144 124 148
rect 144 144 148 148
rect 152 144 156 148
rect 176 144 180 148
rect 120 136 124 140
rect 176 136 180 140
rect 120 128 124 132
rect 176 128 180 132
<< nsubstratencontact >>
rect 132 164 136 168
rect 140 164 144 168
rect 148 164 152 168
rect 156 164 160 168
rect 164 164 168 168
rect 132 156 136 160
rect 164 156 168 160
rect 132 148 136 152
rect 164 148 168 152
rect 132 140 136 144
rect 164 140 168 144
rect 132 132 136 136
rect 164 132 168 136
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_CHAR_c  L500_CHAR_c_0
timestamp 1534321654
transform 1 0 146 0 1 230
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_CHAR_p  L500_CHAR_p_0
timestamp 1534323117
transform 1 0 208 0 1 136
box 0 0 12 18
use L500_CHAR_n  L500_CHAR_n_0
timestamp 1534323210
transform 1 0 224 0 1 136
box 0 0 12 18
use L500_CHAR_p  L500_CHAR_p_1
timestamp 1534323117
transform 1 0 240 0 1 136
box 0 0 12 18
use L500_CHAR_2  L500_CHAR_2_0
timestamp 1534324708
transform 1 0 256 0 1 136
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_CHAR_e  L500_CHAR_e_0
timestamp 1534321786
transform 1 0 114 0 1 50
box 0 0 12 18
use L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 173 0 1 50
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
