magic
tech scmos
timestamp 1541109953
<< error_s >>
rect 3252 2790 3254 3190
rect 3252 1364 3254 1370
rect 3252 1362 3274 1364
rect 3226 1322 3268 1324
rect 3272 1322 3274 1362
rect 3226 1318 3228 1322
rect 3232 1284 3234 1318
rect 3232 1282 3274 1284
rect 3226 1242 3268 1244
rect 3272 1242 3274 1282
rect 3226 1238 3228 1242
rect 3232 1204 3234 1238
rect 3232 1202 3274 1204
rect 3246 1162 3268 1164
rect 3272 1162 3274 1202
rect 3246 1158 3248 1162
rect 3252 1150 3254 1158
rect -226 997 -224 998
rect -227 993 -224 997
rect -227 992 -225 993
rect -227 991 -226 992
rect -175 895 -172 896
rect -118 895 -111 896
rect -103 895 -96 896
rect -174 894 -171 895
rect -173 893 -170 894
rect -172 892 -170 893
rect -95 893 -91 896
rect -86 893 -83 896
rect -43 893 -42 894
rect -95 892 -93 893
rect -85 892 -83 893
rect -44 892 -43 893
rect -171 891 -169 892
rect -45 891 -44 892
rect -171 890 -168 891
rect -46 890 -45 891
rect -171 889 -167 890
rect -47 889 -46 890
rect -169 888 -166 889
rect -168 887 -165 888
rect -51 887 -48 888
rect -167 886 -164 887
rect -51 886 -50 887
rect -167 885 -163 886
rect -52 885 -50 886
rect -165 883 -162 885
rect -54 884 -51 885
rect -55 883 -52 884
rect -163 882 -160 883
rect -56 882 -54 883
rect -162 881 -160 882
rect -57 881 -54 882
rect -161 880 -158 881
rect -59 880 -55 881
rect -160 879 -157 880
rect -61 879 -56 880
rect -396 874 -382 879
rect -159 878 -156 879
rect -62 878 -57 879
rect -158 877 -154 878
rect -157 876 -154 877
rect -64 877 -58 878
rect -64 876 -59 877
rect -155 875 -152 876
rect -66 875 -61 876
rect -154 874 -151 875
rect -67 874 -62 875
rect -445 870 -444 871
rect -406 870 -405 871
rect -446 869 -404 870
rect -445 866 -405 869
rect -445 834 -441 866
rect -435 856 -415 860
rect -435 844 -431 856
rect -419 844 -415 856
rect -435 840 -415 844
rect -409 834 -405 866
rect -445 830 -405 834
rect -391 827 -390 874
rect -387 827 -382 874
rect -152 873 -149 874
rect -104 873 -96 874
rect -69 873 -63 874
rect -151 872 -147 873
rect -106 872 -96 873
rect -71 872 -63 873
rect -150 871 -146 872
rect -148 870 -144 871
rect -107 870 -96 872
rect -72 871 -65 872
rect -73 870 -66 871
rect -147 869 -142 870
rect -107 869 -99 870
rect -96 869 -93 870
rect -74 869 -67 870
rect -76 868 -69 869
rect -114 867 -110 868
rect -101 867 -98 868
rect -76 867 -70 868
rect -101 866 -100 867
rect -79 866 -71 867
rect -80 865 -72 866
rect -81 864 -74 865
rect -82 863 -75 864
rect -84 862 -77 863
rect -84 861 -82 862
rect -86 860 -84 861
rect -391 826 -382 827
rect -448 822 -397 824
rect -448 812 -387 814
rect 663 775 667 776
rect 665 774 666 775
rect 589 762 609 763
rect 585 761 615 762
rect 647 761 649 762
rect 580 760 618 761
rect 646 760 648 761
rect 577 759 591 760
rect 602 759 621 760
rect 645 759 647 760
rect 575 758 587 759
rect 608 758 622 759
rect 644 758 647 759
rect 573 757 583 758
rect 616 757 624 758
rect 643 757 646 758
rect 573 756 582 757
rect 596 756 599 757
rect 601 756 602 757
rect 603 756 605 757
rect 619 756 625 757
rect 642 756 645 757
rect 573 755 580 756
rect 620 755 628 756
rect 640 755 644 756
rect 655 755 657 756
rect 573 754 579 755
rect 621 754 629 755
rect 639 754 643 755
rect 655 754 656 755
rect 568 753 579 754
rect 583 753 584 754
rect 623 753 629 754
rect 638 753 643 754
rect 567 752 579 753
rect 581 752 583 753
rect 566 751 575 752
rect 577 751 583 752
rect 624 752 630 753
rect 638 752 642 753
rect 624 751 631 752
rect 637 751 641 752
rect 565 750 574 751
rect 575 750 580 751
rect 627 750 632 751
rect 565 749 573 750
rect 575 749 579 750
rect 563 748 572 749
rect 575 748 578 749
rect 628 748 633 750
rect 636 749 639 751
rect 563 747 570 748
rect 574 747 576 748
rect 630 747 633 748
rect 562 746 570 747
rect 573 746 576 747
rect 631 746 633 747
rect 634 748 638 749
rect 634 747 637 748
rect 654 747 655 748
rect 634 746 636 747
rect 652 746 655 747
rect 561 745 570 746
rect 572 745 576 746
rect 632 745 636 746
rect 651 745 655 746
rect 560 744 569 745
rect 571 744 575 745
rect 650 744 655 745
rect 560 743 567 744
rect 571 743 573 744
rect 649 743 654 744
rect 557 741 566 743
rect 569 741 572 743
rect 646 742 654 743
rect 646 741 653 742
rect 557 740 564 741
rect 568 740 570 741
rect 555 739 564 740
rect 567 739 570 740
rect 644 740 653 741
rect 658 740 659 741
rect 644 739 651 740
rect 554 738 562 739
rect 553 737 562 738
rect 566 737 568 739
rect 642 738 651 739
rect 656 738 657 739
rect 642 737 649 738
rect 553 736 560 737
rect 563 736 566 737
rect 641 736 647 737
rect 550 735 559 736
rect 563 735 565 736
rect 639 735 647 736
rect 652 735 653 737
rect 549 733 558 735
rect 563 734 564 735
rect 561 733 564 734
rect 547 732 557 733
rect 560 732 563 733
rect 546 731 556 732
rect 559 731 562 732
rect 624 731 625 735
rect 635 734 636 735
rect 639 734 646 735
rect 650 734 652 735
rect 638 733 644 734
rect 634 732 635 733
rect 638 732 643 733
rect 648 732 649 733
rect 633 731 634 732
rect 637 731 642 732
rect 545 730 554 731
rect 559 730 560 731
rect 632 730 634 731
rect 636 730 639 731
rect 545 729 553 730
rect 556 729 559 730
rect 542 728 552 729
rect 555 728 558 729
rect 541 727 551 728
rect 555 727 557 728
rect 540 726 550 727
rect 553 726 556 727
rect 570 726 588 727
rect 624 726 625 730
rect 631 728 633 730
rect 635 729 639 730
rect 634 728 638 729
rect 539 725 550 726
rect 552 725 556 726
rect 569 725 595 726
rect 629 725 632 728
rect 634 727 637 728
rect 634 726 636 727
rect 633 725 636 726
rect 538 724 548 725
rect 551 724 554 725
rect 569 724 599 725
rect 537 723 546 724
rect 551 723 552 724
rect 569 723 574 724
rect 590 723 602 724
rect 536 722 545 723
rect 548 722 551 723
rect 559 722 566 723
rect 534 721 544 722
rect 547 721 550 722
rect 558 721 566 722
rect 532 720 543 721
rect 546 720 549 721
rect 532 719 542 720
rect 545 719 548 720
rect 557 719 566 721
rect 569 722 571 723
rect 594 722 605 723
rect 569 720 570 722
rect 597 721 612 722
rect 578 720 584 721
rect 600 720 614 721
rect 602 719 617 720
rect 530 718 540 719
rect 544 718 546 719
rect 556 718 564 719
rect 566 718 570 719
rect 604 718 620 719
rect 529 717 539 718
rect 543 717 545 718
rect 555 717 562 718
rect 566 717 568 718
rect 607 717 623 718
rect 528 716 537 717
rect 542 716 543 717
rect 554 716 559 717
rect 611 716 623 717
rect 527 715 535 716
rect 540 715 541 716
rect 553 715 558 716
rect 613 715 623 716
rect 624 715 625 725
rect 628 723 636 725
rect 628 721 635 723
rect 631 720 635 721
rect 525 714 533 715
rect 538 714 539 715
rect 552 714 557 715
rect 616 714 623 715
rect 524 713 532 714
rect 551 713 556 714
rect 617 713 623 714
rect 522 712 531 713
rect 536 712 537 713
rect 550 712 554 713
rect 521 711 529 712
rect 549 711 554 712
rect 619 711 623 713
rect 624 711 625 714
rect 630 711 634 719
rect 657 714 672 715
rect 653 713 672 714
rect 636 712 637 713
rect 649 712 669 713
rect 671 712 672 713
rect 520 710 528 711
rect 549 710 553 711
rect 519 709 525 710
rect 548 709 550 710
rect 517 708 523 709
rect 547 708 550 709
rect 635 708 637 712
rect 638 708 641 709
rect 514 707 521 708
rect 512 706 521 707
rect 545 707 549 708
rect 637 707 641 708
rect 545 706 548 707
rect 511 705 518 706
rect 544 705 546 706
rect 510 704 517 705
rect 542 704 546 705
rect 622 704 623 705
rect 508 703 515 704
rect 542 703 545 704
rect 506 702 512 703
rect 541 702 543 703
rect 616 702 623 704
rect 503 701 510 702
rect 540 701 542 702
rect 500 700 508 701
rect 538 700 542 701
rect 616 700 622 702
rect 499 699 507 700
rect 538 699 541 700
rect 616 699 621 700
rect 496 698 505 699
rect 537 698 540 699
rect 616 698 620 699
rect 628 698 629 699
rect 493 697 503 698
rect 536 697 539 698
rect 622 697 629 698
rect 492 696 499 697
rect 536 696 537 697
rect 488 695 497 696
rect 535 695 537 696
rect 487 694 496 695
rect 533 694 536 695
rect 487 693 494 694
rect 532 693 535 694
rect 487 692 492 693
rect 532 692 534 693
rect 487 691 490 692
rect 487 690 489 691
rect 493 690 498 692
rect 531 691 533 692
rect 530 690 533 691
rect 487 689 488 690
rect 493 688 494 690
rect 529 689 531 690
rect 528 688 530 689
rect 528 687 529 688
rect 494 684 495 687
rect 527 686 529 687
rect 526 685 529 686
rect 525 684 529 685
rect 524 683 528 684
rect 524 681 527 683
rect 523 680 526 681
rect 498 678 499 680
rect 522 679 526 680
rect 521 678 526 679
rect 531 678 532 679
rect 521 677 525 678
rect 499 676 501 677
rect 501 675 503 676
rect 520 675 525 677
rect 530 675 531 678
rect 502 674 504 675
rect 520 674 524 675
rect 503 673 507 674
rect 519 673 524 674
rect 504 672 509 673
rect 505 671 511 672
rect 518 671 523 673
rect 525 671 542 675
rect 543 671 555 675
rect 506 670 513 671
rect 518 670 522 671
rect 526 670 528 671
rect 507 669 515 670
rect 517 669 521 670
rect 526 669 527 670
rect 529 669 530 671
rect 542 670 546 671
rect 511 668 516 669
rect 517 668 520 669
rect 541 668 546 670
rect 515 667 519 668
rect 538 667 539 668
rect 540 667 546 668
rect 551 667 552 668
rect 538 666 546 667
rect 550 666 552 667
rect 536 665 545 666
rect 549 665 551 666
rect 535 664 544 665
rect 548 664 550 665
rect 522 661 524 662
rect 535 661 542 664
rect 547 662 548 664
rect 515 659 516 660
rect 515 656 517 659
rect 515 655 518 656
rect 522 655 525 661
rect 532 655 533 661
rect 538 660 542 661
rect 543 660 545 661
rect 543 659 546 660
rect 543 658 547 659
rect 543 657 548 658
rect 544 656 548 657
rect 546 655 549 656
rect 519 652 525 655
rect 538 654 542 655
rect 521 644 525 651
rect 538 648 539 654
rect 540 653 542 654
rect 547 654 550 655
rect 547 653 551 654
rect 563 653 567 654
rect 541 652 542 653
rect 548 651 552 653
rect 564 652 567 653
rect 564 651 566 652
rect 550 650 553 651
rect 551 648 553 650
rect 555 650 560 651
rect 564 650 568 651
rect 555 649 559 650
rect 565 649 568 650
rect 529 644 533 648
rect 538 644 541 648
rect 545 647 547 648
rect 552 647 553 648
rect 554 647 559 649
rect 566 647 568 649
rect 521 641 524 644
rect 540 643 541 644
rect 544 644 547 647
rect 553 646 559 647
rect 554 645 559 646
rect 567 645 569 647
rect 555 644 559 645
rect 544 642 545 644
rect 551 641 556 644
rect 561 643 565 645
rect 560 641 564 643
rect 567 642 570 645
rect 655 644 672 645
rect 654 643 672 644
rect 568 641 570 642
rect 653 642 672 643
rect 653 641 656 642
rect 521 639 523 641
rect 556 640 562 641
rect 563 640 564 641
rect 551 639 555 640
rect 522 638 523 639
rect 522 634 524 638
rect 550 637 555 639
rect 556 637 564 640
rect 569 640 570 641
rect 569 638 572 640
rect 550 636 554 637
rect 559 636 563 637
rect 570 636 572 638
rect 652 638 656 641
rect 660 639 665 642
rect 652 636 655 638
rect 660 637 662 639
rect 549 634 554 636
rect 522 632 525 634
rect 523 630 525 632
rect 549 631 553 634
rect 557 633 559 634
rect 556 631 559 633
rect 523 628 526 630
rect 524 627 526 628
rect 549 629 552 631
rect 555 629 558 631
rect 549 628 551 629
rect 549 627 550 628
rect 555 627 557 629
rect 565 627 567 631
rect 571 630 573 636
rect 652 635 656 636
rect 659 635 662 637
rect 658 634 662 635
rect 573 628 577 630
rect 578 628 581 630
rect 633 629 640 630
rect 633 628 656 629
rect 524 624 527 627
rect 525 622 527 624
rect 569 623 574 627
rect 579 626 580 628
rect 633 627 657 628
rect 579 623 582 626
rect 641 625 647 626
rect 641 623 648 625
rect 569 622 573 623
rect 580 622 583 623
rect 605 622 609 623
rect 641 622 645 623
rect 526 620 528 622
rect 568 620 573 622
rect 581 621 583 622
rect 581 620 584 621
rect 526 618 529 620
rect 567 619 572 620
rect 526 616 530 618
rect 567 617 571 619
rect 566 616 571 617
rect 575 616 579 620
rect 582 617 584 620
rect 606 619 608 622
rect 619 621 626 622
rect 643 621 645 622
rect 619 618 631 621
rect 644 620 646 621
rect 644 619 647 620
rect 654 619 658 627
rect 664 624 665 639
rect 664 619 665 620
rect 644 618 648 619
rect 527 615 531 616
rect 528 613 531 615
rect 566 614 570 616
rect 574 614 576 616
rect 577 615 578 616
rect 583 614 585 617
rect 596 616 601 618
rect 607 617 609 618
rect 645 617 649 618
rect 596 615 600 616
rect 529 612 531 613
rect 529 611 532 612
rect 530 610 532 611
rect 565 611 570 614
rect 573 611 576 614
rect 584 613 586 614
rect 595 613 599 615
rect 608 614 610 617
rect 646 616 649 617
rect 647 615 649 616
rect 661 616 665 619
rect 670 619 671 639
rect 670 616 672 619
rect 661 615 664 616
rect 671 615 672 616
rect 608 613 611 614
rect 584 611 587 613
rect 594 612 599 613
rect 594 611 598 612
rect 530 608 533 610
rect 565 609 569 611
rect 572 609 575 611
rect 585 609 587 611
rect 565 608 568 609
rect 572 608 574 609
rect 531 606 534 608
rect 571 607 574 608
rect 586 607 587 609
rect 593 608 598 611
rect 602 609 606 612
rect 609 611 612 613
rect 610 610 612 611
rect 601 608 605 609
rect 610 608 613 610
rect 532 604 535 606
rect 563 604 567 606
rect 533 603 536 604
rect 534 602 536 603
rect 563 603 566 604
rect 563 602 564 603
rect 571 602 573 607
rect 593 606 597 608
rect 601 607 603 608
rect 611 607 613 608
rect 578 603 581 606
rect 587 604 591 606
rect 588 603 591 604
rect 578 602 580 603
rect 589 602 591 603
rect 534 601 537 602
rect 590 601 591 602
rect 535 599 538 601
rect 588 600 591 601
rect 592 605 597 606
rect 600 605 603 607
rect 612 606 613 607
rect 592 602 596 605
rect 599 602 602 605
rect 612 602 614 606
rect 592 600 595 602
rect 599 600 601 602
rect 613 601 614 602
rect 536 598 539 599
rect 537 597 539 598
rect 590 597 594 600
rect 537 596 540 597
rect 590 596 592 597
rect 598 596 603 600
rect 538 594 541 596
rect 600 594 603 596
rect 605 596 608 600
rect 614 599 618 600
rect 615 597 618 599
rect 616 596 618 597
rect 605 594 606 596
rect 617 594 618 595
rect 628 594 629 615
rect 638 613 643 615
rect 637 611 643 613
rect 648 612 649 615
rect 647 611 649 612
rect 635 609 642 611
rect 646 609 648 611
rect 634 608 640 609
rect 644 608 646 609
rect 634 606 639 608
rect 644 607 645 608
rect 643 606 645 607
rect 649 606 654 607
rect 656 606 660 607
rect 634 605 638 606
rect 640 605 644 606
rect 634 603 637 605
rect 640 603 643 605
rect 649 604 653 606
rect 656 604 659 606
rect 648 603 652 604
rect 656 603 658 604
rect 632 601 635 603
rect 640 602 651 603
rect 656 602 657 603
rect 632 600 634 601
rect 632 599 633 600
rect 539 593 542 594
rect 596 593 603 594
rect 611 593 618 594
rect 540 592 543 593
rect 541 591 544 592
rect 542 590 544 591
rect 619 591 623 594
rect 628 591 631 594
rect 671 591 672 592
rect 619 590 621 591
rect 629 590 631 591
rect 670 590 671 591
rect 543 589 545 590
rect 669 589 670 590
rect 543 588 546 589
rect 668 588 669 589
rect 543 587 547 588
rect 667 587 668 588
rect 545 586 548 587
rect 546 585 549 586
rect 663 585 666 586
rect 547 584 550 585
rect 663 584 664 585
rect 547 583 551 584
rect 662 583 664 584
rect 549 581 552 583
rect 660 582 663 583
rect 659 581 662 582
rect 551 580 554 581
rect 658 580 660 581
rect 552 579 554 580
rect 657 579 660 580
rect 553 578 556 579
rect 655 578 659 579
rect 554 577 557 578
rect 653 577 658 578
rect 555 576 558 577
rect 652 576 657 577
rect 556 575 560 576
rect 557 574 560 575
rect 650 575 656 576
rect 650 574 655 575
rect 559 573 562 574
rect 648 573 653 574
rect 560 572 563 573
rect 647 572 652 573
rect 562 571 565 572
rect 610 571 618 572
rect 645 571 651 572
rect 563 570 567 571
rect 608 570 618 571
rect 643 570 651 571
rect 564 569 568 570
rect 566 568 570 569
rect 607 568 618 570
rect 642 569 649 570
rect 641 568 648 569
rect 567 567 572 568
rect 607 567 615 568
rect 618 567 621 568
rect 640 567 647 568
rect 638 566 645 567
rect 600 565 604 566
rect 613 565 616 566
rect 638 565 644 566
rect 613 564 614 565
rect 635 564 643 565
rect 634 563 642 564
rect 633 562 640 563
rect 632 561 639 562
rect 630 560 637 561
rect 630 559 632 560
rect 628 558 630 559
rect -400 520 -386 525
rect -441 516 -440 517
rect -410 516 -409 517
rect -442 515 -408 516
rect -441 512 -409 515
rect -441 488 -437 512
rect -431 502 -419 506
rect -431 498 -427 502
rect -423 498 -419 502
rect -431 494 -419 498
rect -413 488 -409 512
rect -441 484 -409 488
rect -395 481 -394 520
rect -391 481 -386 520
rect -395 480 -386 481
rect -448 476 -401 478
rect -448 466 -391 468
rect -426 198 -425 200
rect -421 102 -420 198
use contact_meas  contact_meas_0
timestamp 1541109680
transform 1 0 250 0 1 1200
box 0 0 1300 1500
use pnp_table  pnp_table_0
timestamp 1541109953
transform 1 0 -575 0 1 350
box 0 0 300 650
use L500_SIGNATURE_kallisti_big  L500_SIGNATURE_kallisti_big_1 ~/IC/github/PearlRiver/Layout/magic/../../Library/magic
timestamp 1533657739
transform 1 0 -235 0 1 843
box 9 8 231 235
use nmos_table  nmos_table_0
timestamp 1541109953
transform 1 0 750 0 1 850
box 0 0 1700 1700
use metal1_rsquare  metal1_rsquare_0
timestamp 1541109953
transform 0 1 2500 1 0 850
box 0 0 2440 400
use diode_table  diode_table_0
timestamp 1541109953
transform 1 0 50 0 1 850
box 0 0 3104 2800
use metal3_rsquare  metal3_rsquare_0
timestamp 1541109953
transform 0 1 2900 1 0 850
box 0 0 2440 400
use L500_SIGNATURE_kallisti  L500_SIGNATURE_kallisti_0 ~/IC/github/PearlRiver/Layout/magic/../../Library/magic
timestamp 1533657739
transform 1 0 -229 0 1 696
box 4 4 116 118
use L500_SIGNATURE_kallisti  L500_SIGNATURE_kallisti_1
timestamp 1533657739
transform 1 0 -112 0 1 696
box 4 4 116 118
use L500_SIGNATURE_kallisti  L500_SIGNATURE_kallisti_2
timestamp 1533657739
transform 1 0 4 0 1 696
box 4 4 116 118
use hvfet_table  hvfet_table_0
timestamp 1541109953
transform 1 0 -925 0 1 0
box 0 0 650 300
use sonos_table  sonos_table_0
timestamp 1541109953
transform 1 0 -225 0 1 0
box 0 0 650 650
use L500_SIGNATURE_kallisti_big  L500_SIGNATURE_kallisti_big_0
timestamp 1533657739
transform 1 0 479 0 1 541
box 9 8 231 235
use pad_measure  pad_measure_0
timestamp 1541109953
transform 0 1 475 -1 0 504
box 0 0 504 250
use rpoly_rsquare  rpoly_rsquare_0
timestamp 1541109953
transform 1 0 775 0 1 400
box 0 0 2478 400
use ringoscillator_stripe  ringoscillator_stripe_0
timestamp 1541109953
transform 0 1 3360 1 0 450
box 0 0 2704 440
use pmos_table  pmos_table_0
timestamp 1541109953
transform 1 0 3848 0 1 450
box 0 0 1700 1700
use caps_table  caps_table_0
timestamp 1541109953
transform 1 0 3848 0 1 450
box 0 0 2050 2072
use polysi_rsquare  polysi_rsquare_0
timestamp 1541109953
transform 1 0 775 0 1 0
box 0 0 2478 400
use npn_table  npn_table_0
timestamp 1541109953
transform 1 0 3303 0 1 30
box 0 0 650 300
use metal2_rsquare  metal2_rsquare_0
timestamp 1541109953
transform 1 0 4003 0 1 0
box 0 0 2440 400
<< end >>
