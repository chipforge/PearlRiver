magic
tech scmos
timestamp 1531654000
<< nwell >>
rect 0 45 24 64
<< polysilicon >>
rect 7 54 9 56
rect 15 54 17 56
rect 7 44 9 47
rect 3 43 9 44
rect 6 42 9 43
rect 15 44 17 47
rect 15 43 21 44
rect 15 42 18 43
rect 15 29 18 30
rect 15 28 21 29
rect 6 21 9 22
rect 3 20 9 21
rect 7 18 9 20
rect 15 18 17 28
rect 7 8 9 10
rect 15 8 17 10
<< ndiffusion >>
rect 6 10 7 18
rect 9 10 15 18
rect 17 10 18 18
<< pdiffusion >>
rect 2 47 7 54
rect 9 47 15 54
rect 17 47 22 54
<< metal1 >>
rect 0 58 2 62
rect 22 58 24 62
rect 2 47 6 58
rect 10 46 14 54
rect 18 47 22 58
rect 2 30 6 39
rect 2 25 6 26
rect 10 26 14 42
rect 18 38 22 39
rect 18 33 22 34
rect 10 22 22 26
rect 18 18 22 22
rect 2 6 6 10
rect 0 2 2 6
rect 22 2 24 6
<< ntransistor >>
rect 7 10 9 18
rect 15 10 17 18
<< ptransistor >>
rect 7 47 9 54
rect 15 47 17 54
<< polycontact >>
rect 2 39 6 43
rect 18 39 22 43
rect 18 29 22 33
rect 2 21 6 25
<< ndcontact >>
rect 2 10 6 18
rect 18 10 22 18
<< m2contact >>
rect 2 26 6 30
rect 10 42 14 46
rect 18 34 22 38
<< psubstratepcontact >>
rect 2 2 22 6
<< nsubstratencontact >>
rect 2 58 22 62
<< labels >>
rlabel psubstratepcontact 2 2 22 6 1 gnd!
rlabel m2contact 18 34 22 38 7 A
rlabel m2contact 10 42 14 46 1 Z
rlabel m2contact 2 26 6 30 3 B
rlabel nsubstratencontact 2 58 22 62 1 vdd!
<< end >>
