magic
tech scmos
timestamp 1539790345
<< polysilicon >>
rect 130 170 170 186
rect 130 114 170 130
<< metal1 >>
rect 100 226 200 266
rect 100 34 200 74
<< rndiffusion >>
rect 130 154 170 170
<< rpdiffusion >>
rect 130 130 170 146
<< rpoly >>
rect 130 146 170 154
<< polycontact >>
rect 130 186 170 226
rect 130 74 170 114
use L500_TPAD_blank  L500_TPAD_blank_2 ./Library/magic
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
