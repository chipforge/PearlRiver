magic
tech scmos
timestamp 1542691327
<< nwell >>
rect 101 170 199 194
rect 101 130 125 170
rect 175 130 199 170
rect 101 126 132 130
rect 168 126 199 130
rect 101 106 199 126
<< metal1 >>
rect 108 187 192 200
rect 108 170 118 177
rect 182 170 192 177
rect 108 123 118 130
rect 132 134 168 137
rect 182 123 192 130
<< metal2 >>
rect 132 100 168 126
<< nwpbase >>
rect 125 130 175 170
<< pdcontact >>
rect 132 137 168 163
<< m2contact >>
rect 132 126 168 134
<< nsubstratencontact >>
rect 108 177 192 187
rect 108 130 118 170
rect 182 130 192 170
rect 108 113 192 123
use Library/magic/L500_CHAR_d  L500_CHAR_d_0
timestamp 1534321738
transform 1 0 0 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_i  L500_CHAR_i_0
timestamp 1534226087
transform 1 0 16 0 1 304
box 0 0 8 18
use Library/magic/L500_CHAR_o  L500_CHAR_o_1
timestamp 1534323159
transform 1 0 28 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_d  L500_CHAR_d_1
timestamp 1534321738
transform 1 0 44 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_0
timestamp 1534321786
transform 1 0 60 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_under  L500_CHAR_under_0
timestamp 1534325915
transform 1 0 76 0 1 304
box 0 0 12 4
use Library/magic/L500_CHAR_p  L500_CHAR_p_0
timestamp 1534323210
transform 1 0 92 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 108 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_0
timestamp 1534325357
transform 1 0 124 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_s  L500_CHAR_s_1
timestamp 1534323853
transform 1 0 140 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_1
timestamp 1534321786
transform 1 0 156 0 1 304
box 0 0 12 18
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_0
timestamp 1537367970
transform 0 1 0 -1 0 300
box 0 0 100 300
use Library/magic/L500_CHAR_k  L500_CHAR_k_0
timestamp 1534322894
transform 1 0 13 0 1 178
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_2
timestamp 1534325357
transform 1 0 225 0 1 141
box 0 0 12 18
use Library/magic/L500_CHAR_2  L500_CHAR_2_0
timestamp 1534324708
transform 1 0 241 0 1 141
box 0 0 12 18
use Library/magic/L500_CHAR_tick  L500_CHAR_tick_0
timestamp 1541212842
transform 1 0 257 0 1 141
box 0 12 4 18
use Library/magic/L500_CHAR_k  L500_CHAR_k_0
timestamp 1534322894
transform 1 0 265 0 1 141
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_1
timestamp 1534325357
transform 1 0 13 0 1 104
box 0 0 12 18
use Library/magic/L500_METAL2_W100_1rsquare  L500_METAL1_W100_2rsquare_0
timestamp 1537367970
transform 0 1 0 -1 0 100
box 0 0 100 300
<< end >>
