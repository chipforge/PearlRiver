magic
tech scmos
timestamp 1540534681
<< polysilicon >>
rect 140 170 160 188
rect 140 112 160 130
<< metal1 >>
rect 100 226 200 266
rect 140 208 160 226
rect 140 74 160 92
rect 100 34 200 74
<< rndiffusion >>
rect 140 152 160 170
<< rpdiffusion >>
rect 140 130 160 148
<< rpoly >>
rect 140 148 160 152
<< polycontact >>
rect 140 188 160 208
rect 140 92 160 112
use L500_TPAD_blank  L500_TPAD_blank_2 ./Library/magic
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
