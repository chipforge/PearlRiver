magic
tech scmos
timestamp 1534321738
<< metal1 >>
rect 0 17 9 18
rect 0 16 10 17
rect 0 15 11 16
rect 0 14 12 15
rect 0 4 4 14
rect 7 12 12 14
rect 8 6 12 12
rect 7 4 12 6
rect 0 3 12 4
rect 0 2 11 3
rect 0 1 10 2
rect 0 0 9 1
<< end >>
