magic
tech scmos
timestamp 1540533394
<< polysilicon >>
rect 147 165 152 171
rect 147 130 152 136
<< metal1 >>
rect 90 181 100 200
rect 200 181 210 200
rect 90 171 145 181
rect 155 171 210 181
rect 90 120 145 130
rect 155 120 210 130
rect 90 100 100 120
rect 200 100 210 120
<< rndiffusion >>
rect 147 153 152 159
<< rpdiffusion >>
rect 147 142 152 148
<< rpoly >>
rect 147 148 152 153
<< polycontact >>
rect 145 171 155 181
rect 145 120 155 130
<< polyndiff >>
rect 147 159 152 165
<< polypdiff >>
rect 147 136 152 142
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
