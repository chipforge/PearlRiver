magic
tech scmos
timestamp 1534324785
<< metal1 >>
rect 0 17 10 18
rect 0 16 11 17
rect 0 14 12 16
rect 6 13 12 14
rect 8 10 12 13
rect 0 7 12 10
rect 8 4 12 7
rect 6 3 12 4
rect 0 2 12 3
rect 0 1 11 2
rect 0 0 10 1
<< end >>
