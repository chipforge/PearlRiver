magic
tech scmos
timestamp 1539788087
<< polysilicon >>
rect 130 160 170 168
rect 130 132 170 140
<< metal1 >>
rect 100 208 210 248
rect 100 52 200 92
<< rndiffusion >>
rect 130 152 170 160
<< rpdiffusion >>
rect 130 140 170 148
<< rpoly >>
rect 130 148 170 152
<< polycontact >>
rect 130 168 170 208
rect 130 92 170 132
use L500_TPAD_blank  L500_TPAD_blank_1 ./Library/magic
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
