magic
tech scmos
timestamp 1539785150
<< polysilicon >>
rect 130 157 170 163
rect 130 137 170 143
<< metal1 >>
rect 100 203 200 243
rect 100 57 200 97
<< rndiffusion >>
rect 130 151 170 157
<< rpdiffusion >>
rect 130 143 170 149
<< rpoly >>
rect 130 149 170 151
<< polycontact >>
rect 130 163 170 203
rect 130 97 170 137
use L500_TPAD_blank  L500_TPAD_blank_1 ./Library/magic
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
