magic
tech scmos
timestamp 1533885931
<< metal2 >>
rect 1170 468 1174 470
rect 2434 446 2438 448
rect 2042 300 2046 302
rect 378 294 382 296
rect 378 188 382 190
rect 1170 -2 1174 0
use Library/magic/L500_TPM2_blank  L500_TPM2_blank_2 Library/magic
timestamp 1533879882
transform 1 0 1072 0 1 462
box 0 0 120 120
use Library/magic/L500_TPM2_blank  L500_TPM2_blank_4
timestamp 1533879882
transform 1 0 2336 0 1 440
box 0 0 120 120
use Layout/magic/T7_RO51_INV  T7_RO51_INV_0 Layout/magic
timestamp 1533818910
transform 1 0 2024 0 1 310
box -360 -8 784 136
use Layout/magic/T10_RO51_NAND3  T10_RO51_NAND3_0
timestamp 1533837380
transform 1 0 360 0 1 304
box -360 -8 1184 164
use Library/magic/L500_TPM2_blank  L500_TPM2_blank_3
timestamp 1533879882
transform 1 0 1944 0 1 188
box 0 0 120 120
use Library/magic/L500_TPM2_blank  L500_TPM2_blank_0
timestamp 1533879882
transform 1 0 360 0 1 182
box 0 0 120 120
use Layout/magic/T7_CELL50_FILLCAP  T7_CELL50_FILLCAP_0
timestamp 1533830913
transform 1 0 2024 0 1 40
box -360 -2 960 130
use Layout/magic/T11_RO51_NOR3  T11_RO51_NOR3_0
timestamp 1533837380
transform 1 0 360 0 -1 180
box -360 -8 1184 180
use Library/magic/L500_TPM2_blank  L500_TPM2_blank_1
timestamp 1533879882
transform 1 0 1072 0 1 -114
box 0 0 120 120
<< end >>
