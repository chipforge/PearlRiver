magic
tech scmos
timestamp 1531674175
<< nwell >>
rect 0 32 24 48
<< polysilicon >>
rect 7 38 9 40
rect 15 38 17 40
rect 7 32 9 35
rect 3 31 9 32
rect 6 30 9 31
rect 15 32 17 35
rect 15 31 21 32
rect 15 30 18 31
rect 6 17 9 18
rect 3 16 9 17
rect 7 13 9 16
rect 15 17 18 18
rect 15 16 21 17
rect 15 13 17 16
rect 7 8 9 10
rect 15 8 17 10
<< ndiffusion >>
rect 6 10 7 13
rect 9 10 15 13
rect 17 10 18 13
<< pdiffusion >>
rect 6 35 7 38
rect 9 35 10 38
rect 14 35 15 38
rect 17 35 18 38
<< metal1 >>
rect 0 42 2 46
rect 22 42 24 46
rect 2 38 6 42
rect 18 38 22 42
rect 2 26 6 27
rect 2 21 6 22
rect 10 26 14 34
rect 10 14 14 22
rect 18 26 22 27
rect 18 21 22 22
rect 10 10 18 14
rect 2 6 6 10
rect 0 2 2 6
rect 22 2 24 6
<< ntransistor >>
rect 7 10 9 13
rect 15 10 17 13
<< ptransistor >>
rect 7 35 9 38
rect 15 35 17 38
<< polycontact >>
rect 2 27 6 31
rect 18 27 22 31
rect 2 17 6 21
rect 18 17 22 21
<< ndcontact >>
rect 2 10 6 14
rect 18 10 22 14
<< pdcontact >>
rect 2 34 6 38
rect 10 34 14 38
rect 18 34 22 38
<< m2contact >>
rect 2 22 6 26
rect 10 22 14 26
rect 18 22 22 26
<< psubstratepcontact >>
rect 2 2 22 6
<< nsubstratencontact >>
rect 2 42 22 46
<< labels >>
rlabel psubstratepcontact 2 2 22 6 1 gnd!
rlabel m2contact 18 22 22 26 1 A
rlabel m2contact 2 22 6 26 3 B
rlabel m2contact 10 22 14 26 1 Z
rlabel nsubstratencontact 2 42 22 46 5 vdd!
<< end >>
