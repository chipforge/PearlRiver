magic
tech scmos
timestamp 1540534609
<< polysilicon >>
rect 140 158 160 165
rect 140 136 160 143
<< metal1 >>
rect 100 203 200 223
rect 140 185 160 203
rect 140 97 160 116
rect 100 77 200 97
<< rndiffusion >>
rect 140 151 160 158
<< rpdiffusion >>
rect 140 143 160 150
<< rpoly >>
rect 140 150 160 151
<< polycontact >>
rect 140 165 160 185
rect 140 116 160 136
use L500_TPAD_blank  L500_TPAD_blank_1 ./Library/magic
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
