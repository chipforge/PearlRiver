magic
tech scmos
timestamp 1540534869
<< polysilicon >>
rect 145 160 155 169
rect 145 131 155 140
<< metal1 >>
rect 100 200 200 210
rect 145 179 155 200
rect 145 100 155 121
rect 100 90 200 100
<< rndiffusion >>
rect 145 151 155 160
<< rpdiffusion >>
rect 145 140 155 149
<< rpoly >>
rect 145 149 155 151
<< polycontact >>
rect 145 169 155 179
rect 145 121 155 131
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
