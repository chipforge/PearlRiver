magic
tech scmos
timestamp 1531585550
<< nwell >>
rect 0 56 32 88
<< polysilicon >>
rect 7 78 9 80
rect 15 78 17 80
rect 23 78 25 80
rect 7 56 9 58
rect 3 55 9 56
rect 6 54 9 55
rect 15 52 17 58
rect 11 51 17 52
rect 14 50 17 51
rect 23 48 25 58
rect 19 47 25 48
rect 22 46 25 47
rect 22 25 25 26
rect 11 22 13 25
rect 19 24 25 25
rect 11 20 17 22
rect 6 17 9 18
rect 3 16 9 17
rect 7 14 9 16
rect 15 14 17 20
rect 23 14 25 24
rect 7 8 9 10
rect 15 8 17 10
rect 23 8 25 10
<< ndiffusion >>
rect 6 10 7 14
rect 9 10 10 14
rect 14 10 15 14
rect 17 10 18 14
rect 22 10 23 14
rect 25 10 26 14
<< pdiffusion >>
rect 6 58 7 78
rect 9 58 15 78
rect 17 58 23 78
rect 25 58 26 78
<< metal1 >>
rect 0 82 2 86
rect 30 82 32 86
rect 2 78 6 82
rect 26 54 30 58
rect 2 30 6 51
rect 2 21 6 26
rect 10 46 14 47
rect 10 29 14 42
rect 18 38 22 43
rect 18 29 22 34
rect 26 22 30 50
rect 10 18 30 22
rect 10 14 14 18
rect 26 14 30 18
rect 2 6 6 10
rect 18 6 22 10
rect 0 2 2 6
rect 30 2 32 6
<< ntransistor >>
rect 7 10 9 14
rect 15 10 17 14
rect 23 10 25 14
<< ptransistor >>
rect 7 58 9 78
rect 15 58 17 78
rect 23 58 25 78
<< polycontact >>
rect 2 51 6 55
rect 10 47 14 51
rect 18 43 22 47
rect 10 25 14 29
rect 18 25 22 29
rect 2 17 6 21
<< ndcontact >>
rect 2 10 6 14
rect 10 10 14 14
rect 18 10 22 14
rect 26 10 30 14
<< pdcontact >>
rect 2 58 6 78
rect 26 58 30 78
<< m2contact >>
rect 2 82 30 86
rect 2 26 6 30
rect 26 50 30 54
rect 10 42 14 46
rect 18 34 22 38
rect 2 2 30 6
<< psubstratepcontact >>
rect 0 2 30 6
<< nsubstratencontact >>
rect 0 82 30 86
<< labels >>
rlabel nsubstratencontact 2 82 30 86 5 vdd!
rlabel psubstratepcontact 2 2 30 6 1 gnd!
rlabel m2contact 18 34 22 38 1 A
rlabel m2contact 26 50 30 54 1 Z
rlabel m2contact 10 42 14 46 1 B
rlabel m2contact 2 26 6 30 3 C
<< end >>
