magic
tech scmos
timestamp 1540534943
<< polysilicon >>
rect 145 166 155 181
rect 145 118 155 133
<< metal1 >>
rect 90 191 100 200
rect 200 191 210 200
rect 90 181 145 191
rect 155 181 210 191
rect 90 108 145 118
rect 155 108 210 118
rect 90 100 100 108
rect 200 100 210 108
<< rndiffusion >>
rect 145 151 155 166
<< rpdiffusion >>
rect 145 133 155 148
<< rpoly >>
rect 145 148 155 151
<< polycontact >>
rect 145 181 155 191
rect 145 108 155 118
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
