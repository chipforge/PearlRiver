magic
tech scmos
timestamp 1531599168
use Library/magic/T10_NAND3  T10_NAND3_49 Library/magic
timestamp 1531593415
transform -1 0 32 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_48
timestamp 1531593415
transform -1 0 64 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_47
timestamp 1531593415
transform -1 0 96 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_46
timestamp 1531593415
transform -1 0 128 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_45
timestamp 1531593415
transform -1 0 160 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_44
timestamp 1531593415
transform -1 0 192 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_43
timestamp 1531593415
transform -1 0 224 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_42
timestamp 1531593415
transform -1 0 256 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_41
timestamp 1531593415
transform -1 0 288 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_40
timestamp 1531593415
transform -1 0 320 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_39
timestamp 1531593415
transform -1 0 352 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_38
timestamp 1531593415
transform -1 0 384 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_37
timestamp 1531593415
transform -1 0 416 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_36
timestamp 1531593415
transform -1 0 448 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_35
timestamp 1531593415
transform -1 0 480 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_34
timestamp 1531593415
transform -1 0 512 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_33
timestamp 1531593415
transform -1 0 544 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_32
timestamp 1531593415
transform -1 0 576 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_31
timestamp 1531593415
transform -1 0 608 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_30
timestamp 1531593415
transform -1 0 640 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_29
timestamp 1531593415
transform -1 0 672 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_28
timestamp 1531593415
transform -1 0 704 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_27
timestamp 1531593415
transform -1 0 736 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_26
timestamp 1531593415
transform -1 0 768 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_25
timestamp 1531593415
transform -1 0 800 0 -1 158
box 0 2 32 80
use Library/magic/T10_NAND2  T10_NAND2_1 Library/magic
timestamp 1531593307
transform -1 0 824 0 -1 158
box 0 2 24 80
use Library/magic/T10_NAND2  T10_NAND2_0
timestamp 1531593307
transform 1 0 0 0 1 -2
box 0 2 24 80
use Library/magic/T10_NAND3  T10_NAND3_0
timestamp 1531593415
transform 1 0 24 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_1
timestamp 1531593415
transform 1 0 56 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_2
timestamp 1531593415
transform 1 0 88 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_3
timestamp 1531593415
transform 1 0 120 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_4
timestamp 1531593415
transform 1 0 152 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_5
timestamp 1531593415
transform 1 0 184 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_6
timestamp 1531593415
transform 1 0 216 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_7
timestamp 1531593415
transform 1 0 248 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_8
timestamp 1531593415
transform 1 0 280 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_9
timestamp 1531593415
transform 1 0 312 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_10
timestamp 1531593415
transform 1 0 344 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_11
timestamp 1531593415
transform 1 0 376 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_12
timestamp 1531593415
transform 1 0 408 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_13
timestamp 1531593415
transform 1 0 440 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_14
timestamp 1531593415
transform 1 0 472 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_15
timestamp 1531593415
transform 1 0 504 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_16
timestamp 1531593415
transform 1 0 536 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_17
timestamp 1531593415
transform 1 0 568 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_18
timestamp 1531593415
transform 1 0 600 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_19
timestamp 1531593415
transform 1 0 632 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_20
timestamp 1531593415
transform 1 0 664 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_21
timestamp 1531593415
transform 1 0 696 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_22
timestamp 1531593415
transform 1 0 728 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_23
timestamp 1531593415
transform 1 0 760 0 1 -2
box 0 2 32 80
use Library/magic/T10_NAND3  T10_NAND3_24
timestamp 1531593415
transform 1 0 792 0 1 -2
box 0 2 32 80
<< end >>
