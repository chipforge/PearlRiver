magic
tech scmos
timestamp 1534323034
<< metal1 >>
rect 2 17 5 18
rect 11 17 14 18
rect 1 16 6 17
rect 10 16 15 17
rect 0 12 16 16
rect 0 0 4 12
rect 7 0 10 12
rect 13 0 16 12
<< end >>
