magic
tech scmos
timestamp 1538237708
use Library/magic/L500_METAL1_W4m_100rsquare  L500_METAL1_W4m_100rsquare_0 Library/magic
timestamp 1537372519
transform 1 0 200 0 1 300
box 0 0 420 100
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_4 Library/magic
timestamp 1537367970
transform 0 1 520 -1 0 400
box 0 0 100 300
use Library/magic/L500_METAL1_W4_100rsquare  L500_METAL1_W4_100rsquare_0 Library/magic
timestamp 1537368500
transform 1 0 1840 0 1 300
box 0 0 600 100
use Library/magic/L500_METAL1_W10_100rsquare  L500_METAL1_W10_100rsquare_0 Library/magic
timestamp 1537368500
transform 1 0 0 0 1 200
box 0 0 1200 100
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_1
timestamp 1537367970
transform 0 1 1100 -1 0 300
box 0 0 100 300
use Library/magic/L500_METAL1_W6_100rsquare  L500_METAL1_W6_100rsquare_0 Library/magic
timestamp 1537368500
transform 1 0 1300 0 1 200
box 0 0 800 100
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_2
timestamp 1537367970
transform 0 1 2000 -1 0 300
box 0 0 100 300
use Library/magic/L500_METAL2_W100_1rsquare  L500_METAL2_W100_1rsquare_0 Library/magic
timestamp 1537367970
transform 1 0 200 0 1 100
box 0 0 100 300
use Library/magic/L500_METAL1_W8m_100rsquare  L500_METAL1_W8m_100rsquare_0 Library/magic
timestamp 1537373212
transform 1 0 200 0 1 100
box 0 0 640 100
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_5
timestamp 1537367970
transform 0 1 740 -1 0 200
box 0 0 100 300
use Library/magic/L500_METAL1_W8_100rsquare  L500_METAL1_W8_100rsquare_0 Library/magic
timestamp 1537368500
transform 1 0 940 0 1 100
box 0 0 1000 100
use Library/magic/L500_METAL2_W100_1rsquare  L500_METAL2_W100_1rsquare_1
timestamp 1537367970
transform -1 0 1940 0 -1 400
box 0 0 100 300
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_6
timestamp 1537367970
transform 1 0 2340 0 1 100
box 0 0 100 300
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_0
timestamp 1537367970
transform 1 0 0 0 1 0
box 0 0 100 300
use Library/magic/L500_METAL1_W19_100rsquare  L500_METAL1_190_100rsquare_0 Library/magic
timestamp 1537368500
transform 1 0 0 0 1 0
box 0 0 2100 100
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_3
timestamp 1537367970
transform 0 1 2000 -1 0 100
box 0 0 100 300
<< end >>
