magic
tech scmos
timestamp 1534327497
<< metal1 >>
rect 2 17 10 18
rect 1 16 11 17
rect 0 14 12 16
rect 0 10 4 14
rect 8 10 12 14
rect 0 8 12 10
rect 1 7 12 8
rect 2 6 12 7
rect 8 3 12 6
rect 0 2 12 3
rect 0 0 11 2
<< end >>
