magic
tech scmos
timestamp 1538471569
<< nwell >>
rect 6 5 60 34
<< metal1 >>
rect 14 5 19 17
rect 31 5 36 17
rect 45 5 50 17
<< collector >>
rect 12 22 21 24
rect 12 17 14 22
rect 19 17 21 22
rect 12 15 21 17
<< emitter >>
rect 29 22 38 24
rect 29 17 31 22
rect 36 17 38 22
rect 29 15 38 17
<< pbase >>
rect 25 24 54 28
rect 25 15 29 24
rect 38 22 54 24
rect 38 17 45 22
rect 50 17 54 22
rect 38 15 54 17
rect 25 11 54 15
<< collectorcontact >>
rect 14 17 19 22
<< emittercontact >>
rect 31 17 36 22
<< pbasecontact >>
rect 45 17 50 22
<< end >>
