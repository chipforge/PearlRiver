magic
tech scmos
timestamp 1540543464
<< polysilicon >>
rect 145 166 155 181
rect 145 118 155 133
<< metal1 >>
rect 90 191 100 200
rect 200 191 210 200
rect 90 181 145 191
rect 155 181 210 191
rect 90 108 145 118
rect 155 108 210 118
rect 90 100 100 108
rect 200 100 210 108
<< rndiffusion >>
rect 145 151 155 166
<< rpdiffusion >>
rect 145 133 155 148
<< rpoly >>
rect 145 148 155 151
<< polycontact >>
rect 145 181 155 191
rect 145 108 155 118
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use Library/magic/L500_CHAR_k  L500_CHAR_k_0
timestamp 1534322894
transform 1 0 145 0 1 220
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use Library/magic/L500_CHAR_d  L500_CHAR_d_0
timestamp 1534321738
transform 1 0 225 0 1 140
box 0 0 12 18
use Library/magic/L500_CHAR_w  L500_CHAR_w_0
timestamp 1534324213
transform 1 0 244 0 1 151
box 0 0 16 18
use Library/magic/L500_CHAR_1  L500_CHAR_1_0
timestamp 1534326485
transform 1 0 264 0 1 151
box 0 0 12 18
use Library/magic/L500_CHAR_0  L500_CHAR_0_0
timestamp 1534325425
transform 1 0 280 0 1 151
box 0 0 12 18
use Library/magic/L500_CHAR_slash  L500_CHAR_slash_0
timestamp 1534532558
transform 1 0 296 0 1 151
box 0 0 8 18
use Library/magic/L500_CHAR_l  L500_CHAR_l_0
timestamp 1534225390
transform 1 0 244 0 1 129
box 0 0 12 18
use Library/magic/L500_CHAR_3  L500_CHAR_3_1
timestamp 1534324785
transform 1 0 260 0 1 129
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use Library/magic/L500_CHAR_a  L500_CHAR_a_0
timestamp 1534325357
transform 1 0 145 0 1 60
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
