magic
tech scmos
timestamp 1539785774
<< polysilicon >>
rect 140 160 160 168
rect 140 132 160 140
<< metal1 >>
rect 100 200 200 220
rect 140 188 160 200
rect 140 100 160 112
rect 100 80 200 100
<< rndiffusion >>
rect 140 152 160 160
<< rpdiffusion >>
rect 140 140 160 148
<< rpoly >>
rect 140 148 160 152
<< polycontact >>
rect 140 168 160 188
rect 140 112 160 132
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
