magic
tech scmos
timestamp 1534224731
<< metal1 >>
rect 0 10 4 18
rect 8 10 12 18
rect 0 6 12 10
rect 0 0 4 6
rect 8 0 12 6
<< end >>
