magic
tech scmos
timestamp 1541105680
<< error_s >>
rect 175 170 189 175
rect 134 166 135 167
rect 165 166 166 167
rect 133 165 167 166
rect 134 162 166 165
rect 134 138 138 162
rect 144 152 156 156
rect 144 148 148 152
rect 152 148 156 152
rect 144 144 156 148
rect 162 138 166 162
rect 134 134 166 138
rect 180 131 181 170
rect 184 131 189 170
rect 180 130 189 131
rect 126 126 174 128
rect 116 116 184 118
<< nwell >>
rect 110 174 190 190
rect 110 126 126 174
rect 138 156 162 162
rect 138 144 144 156
rect 156 144 162 156
rect 138 138 162 144
rect 174 126 190 174
rect 110 118 190 126
<< metal1 >>
rect 100 208 200 218
rect 145 172 155 208
rect 128 170 172 172
rect 128 130 130 170
rect 134 164 166 166
rect 134 130 136 164
rect 128 128 136 130
rect 146 85 154 154
rect 164 130 166 164
rect 170 130 172 170
rect 164 128 172 130
rect 178 170 186 172
rect 178 130 180 170
rect 184 130 186 170
rect 100 75 154 85
rect 178 90 186 130
rect 178 80 200 90
<< nwpbase >>
rect 126 162 174 174
rect 126 138 138 162
rect 144 144 156 156
rect 162 138 174 162
rect 126 126 174 138
<< pbasepdiffcontact >>
rect 148 148 152 152
<< ndcontact >>
rect 180 130 184 170
<< pdcontact >>
rect 130 166 170 170
rect 130 130 134 166
rect 166 130 170 166
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_CHAR_c  L500_CHAR_c_0
timestamp 1534321654
transform 1 0 146 0 1 230
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_CHAR_p  L500_CHAR_p_0
timestamp 1534323210
transform 1 0 208 0 1 136
box 0 0 12 18
use L500_CHAR_n  L500_CHAR_n_0
timestamp 1534323117
transform 1 0 224 0 1 136
box 0 0 12 18
use L500_CHAR_p  L500_CHAR_p_1
timestamp 1534323210
transform 1 0 240 0 1 136
box 0 0 12 18
use L500_CHAR_1  L500_CHAR_1_0
timestamp 1534326485
transform 1 0 256 0 1 136
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_CHAR_e  L500_CHAR_e_0
timestamp 1534321786
transform 1 0 114 0 1 50
box 0 0 12 18
use L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 173 0 1 50
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
