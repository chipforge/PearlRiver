magic
tech scmos
timestamp 1541236225
<< nwell >>
rect 26 175 274 199
rect 26 125 50 175
rect 250 125 274 175
rect 26 121 57 125
rect 107 121 274 125
rect 26 101 274 121
<< metal1 >>
rect 33 192 267 200
rect 33 175 43 182
rect 257 175 267 182
rect 33 118 43 125
rect 57 129 243 168
rect 257 118 267 125
<< metal2 >>
rect 57 100 243 121
<< nwpbase >>
rect 50 125 250 175
rect 57 121 107 125
<< pbasendiffcontact >>
rect 57 132 243 168
<< m2contact >>
rect 57 121 243 129
<< nsubstratencontact >>
rect 33 182 267 192
rect 33 125 43 175
rect 257 125 267 175
rect 33 108 267 118
use Library/magic/L500_CHAR_d  L500_CHAR_d_0
timestamp 1534321738
transform 1 0 0 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_i  L500_CHAR_i_0
timestamp 1534226087
transform 1 0 16 0 1 304
box 0 0 8 18
use Library/magic/L500_CHAR_o  L500_CHAR_o_1
timestamp 1534323159
transform 1 0 28 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_d  L500_CHAR_d_1
timestamp 1534321738
transform 1 0 44 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_0
timestamp 1534321786
transform 1 0 60 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_under  L500_CHAR_under_0
timestamp 1534325915
transform 1 0 76 0 1 304
box 0 0 12 4
use Library/magic/L500_CHAR_p  L500_CHAR_p_0
timestamp 1534323210
transform 1 0 92 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 108 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_0
timestamp 1534325357
transform 1 0 124 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_s  L500_CHAR_s_1
timestamp 1534323853
transform 1 0 140 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_1
timestamp 1534321786
transform 1 0 156 0 1 304
box 0 0 12 18
use Library/magic/L500_METAL1_W100_1rsquare  L500_METAL1_W100_1rsquare_0
timestamp 1537367970
transform 0 1 0 -1 0 300
box 0 0 100 300
use Library/magic/L500_CHAR_k  L500_CHAR_k_0
timestamp 1534322894
transform 1 0 13 0 1 178
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_2
timestamp 1534325357
transform 1 0 273 0 1 163
box 0 0 12 18
use Library/magic/L500_CHAR_1  L500_CHAR_1_0
timestamp 1534326485
transform 1 0 273 0 1 141
box 0 0 12 18
use Library/magic/L500_CHAR_0  L500_CHAR_0_1
timestamp 1534325425
transform 1 0 289 0 1 141
box 0 0 12 18
use Library/magic/L500_CHAR_tick  L500_CHAR_tick_0
timestamp 1541212842
transform 1 0 273 0 1 119
box 0 12 4 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_1
timestamp 1534325357
transform 1 0 13 0 1 104
box 0 0 12 18
use Library/magic/L500_CHAR_k  Library/magic/L500_CHAR_k_0
timestamp 1534322894
transform 1 0 281 0 1 119
box 0 0 12 18
use Library/magic/L500_METAL2_W100_1rsquare  L500_METAL1_W100_2rsquare_0
timestamp 1537367970
transform 0 1 0 -1 0 100
box 0 0 100 300
<< end >>
