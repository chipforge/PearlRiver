magic
tech scmos
timestamp 1542092493
<< error_s >>
rect 148 151 151 152
use Library/magic/L500_NMOSi_W40_L40_params  L500_NMOSi_W40_L40_params_0
timestamp 1542090445
transform 1 0 0 0 1 1400
box 0 0 300 300
use Library/magic/L500_NMOSi_W20_L20_params  L500_NMOSi_W20_L20_params_0
timestamp 1542090445
transform 1 0 0 0 1 1050
box 0 0 300 300
use Library/magic/L500_NMOSi_W10_L10_params  L500_NMOSi_W10_L10_params_0
timestamp 1542090445
transform 1 0 0 0 1 700
box 0 0 300 300
use Library/magic/L500_NMOSi_W5_L5_params  L500_NMOSi_W5_L5_params_0
timestamp 1542090445
transform 1 0 0 0 1 350
box 0 0 300 300
use Library/magic/L500_NMOSi_W3_L2_params  L500_NMOSi_W3_L2_params_0
timestamp 1542090651
transform 1 0 0 0 1 0
box 0 0 300 300
<< end >>
