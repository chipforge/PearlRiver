magic
tech scmos
timestamp 1534323210
<< metal1 >>
rect 2 17 10 18
rect 1 16 11 17
rect 0 14 12 16
rect 0 10 4 14
rect 8 11 12 14
rect 7 10 12 11
rect 0 9 12 10
rect 0 8 11 9
rect 0 7 10 8
rect 0 6 9 7
rect 0 0 4 6
<< end >>
