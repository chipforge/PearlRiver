magic
tech scmos
timestamp 1540535036
<< polysilicon >>
rect 145 165 155 178
rect 145 122 155 135
<< metal1 >>
rect 90 188 100 200
rect 200 188 210 200
rect 90 178 145 188
rect 155 178 210 188
rect 90 112 145 122
rect 155 112 210 122
rect 90 100 100 112
rect 200 100 210 112
<< rndiffusion >>
rect 145 152 155 165
<< rpdiffusion >>
rect 145 135 155 148
<< rpoly >>
rect 145 148 155 152
<< polycontact >>
rect 145 178 155 188
rect 145 112 155 122
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
