magic
tech scmos
timestamp 1538326853
<< polysilicon >>
rect 107 48 503 52
<< metal1 >>
rect 100 48 103 52
rect 507 48 510 52
<< polycontact >>
rect 103 48 107 52
rect 503 48 507 52
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_1 Library/magic
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 510 0 1 0
box 0 0 100 100
<< end >>
