magic
tech scmos
timestamp 1534324213
<< metal1 >>
rect 0 5 4 18
rect 7 5 10 18
rect 13 5 16 18
rect 0 2 16 5
rect 1 1 7 2
rect 10 1 15 2
rect 2 0 5 1
rect 11 0 14 1
<< end >>
