magic
tech scmos
timestamp 1534321816
<< metal1 >>
rect 2 16 12 18
rect 0 14 12 16
rect 0 10 4 14
rect 0 6 10 10
rect 0 0 4 6
<< end >>
