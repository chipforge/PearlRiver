magic
tech scmos
timestamp 1534226087
<< metal1 >>
rect 0 14 8 18
rect 2 4 6 14
rect 0 0 8 4
<< end >>
