magic
tech scmos
timestamp 1531593307
<< nwell >>
rect 0 60 24 80
<< polysilicon >>
rect 7 70 9 72
rect 15 70 17 72
rect 7 60 9 62
rect 3 59 9 60
rect 6 58 9 59
rect 15 60 17 62
rect 15 59 21 60
rect 15 58 18 59
rect 15 29 18 30
rect 15 28 21 29
rect 6 21 9 22
rect 3 20 9 21
rect 7 18 9 20
rect 15 18 17 28
rect 7 8 9 10
rect 15 8 17 10
<< ndiffusion >>
rect 6 10 7 18
rect 9 10 15 18
rect 17 10 18 18
<< pdiffusion >>
rect 6 62 7 70
rect 9 62 10 70
rect 14 62 15 70
rect 17 62 18 70
<< metal1 >>
rect 0 74 2 78
rect 22 74 24 78
rect 2 70 6 74
rect 18 70 22 74
rect 2 46 6 55
rect 2 25 6 42
rect 10 54 14 62
rect 10 26 14 50
rect 18 38 22 55
rect 18 33 22 34
rect 10 22 22 26
rect 18 18 22 22
rect 2 6 6 10
rect 0 2 2 6
rect 22 2 24 6
<< ntransistor >>
rect 7 10 9 18
rect 15 10 17 18
<< ptransistor >>
rect 7 62 9 70
rect 15 62 17 70
<< polycontact >>
rect 2 55 6 59
rect 18 55 22 59
rect 18 29 22 33
rect 2 21 6 25
<< ndcontact >>
rect 2 10 6 18
rect 18 10 22 18
<< pdcontact >>
rect 2 62 6 70
rect 10 62 14 70
rect 18 62 22 70
<< m2contact >>
rect 2 42 6 46
rect 10 50 14 54
rect 18 34 22 38
<< psubstratepcontact >>
rect 2 2 22 6
<< nsubstratencontact >>
rect 2 74 22 78
<< labels >>
rlabel psubstratepcontact 2 2 22 6 1 gnd!
rlabel nsubstratencontact 2 74 22 78 5 vdd!
rlabel m2contact 18 34 22 38 7 A
rlabel m2contact 10 50 14 54 1 Z
rlabel m2contact 2 42 6 46 3 B
<< end >>
