magic
tech scmos
timestamp 1540677881
<< error_p >>
rect -30 92 -17 97
rect -15 92 -4 97
rect -22 -7 -17 92
rect -30 -8 -17 -7
rect -10 -7 -9 92
rect -4 -7 1 92
rect -10 -8 1 -7
<< nwell >>
rect -48 104 70 116
rect -48 -20 -4 104
rect 58 -20 70 104
rect -48 -32 70 -20
<< polysilicon >>
rect -16 92 6 96
rect -16 -8 -10 92
rect -16 -12 6 -8
<< ndiffusion >>
rect -36 90 -22 92
rect -36 -6 -34 90
rect -24 -6 -22 90
rect -36 -8 -22 -6
<< metal1 >>
rect -36 90 -22 92
rect -36 -6 -34 90
rect -24 -6 -22 90
rect -36 -8 -22 -6
rect 6 90 46 92
rect 6 -6 10 90
rect 20 -6 34 90
rect 44 -6 46 90
rect 6 -8 46 -6
<< ntransistor >>
rect -10 -8 6 92
<< nwpbase >>
rect -4 -20 58 104
<< pbasendiffusion >>
rect 6 90 22 92
rect 6 -6 10 90
rect 20 -6 22 90
rect 6 -8 22 -6
<< pbasepdiffusion >>
rect 32 90 46 92
rect 32 -6 34 90
rect 44 -6 46 90
rect 32 -8 46 -6
<< ndcontact >>
rect -34 -6 -24 90
rect 10 -6 20 90
<< pdcontact >>
rect 34 -6 44 90
<< end >>
